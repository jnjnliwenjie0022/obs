`ifdef ATCBMC300_CONST_VH
`else
`define ATCBMC300_CONST_VH
`define ATCBMC300_PRODUCT_ID 32'h00003005

`define ATCBMC300_SLV0_SIZE 1
//VPERL_BEGIN
//	for($i=0;$i<16;$i++) {
//		for($j=0;$j<32;$j++) {
// :`ifdef ATCBMC300_MST${i}_SLV${j} 
// :	`define ATCBMC300_M${i}S${j} 1'b1 
// :`else 
// :	`define ATCBMC300_M${i}S${j} 1'b0 
// :`endif 
//		}
//	}
//VPERL_END

// VPERL_GENERATED_BEGIN
`ifdef ATCBMC300_MST0_SLV0
	`define ATCBMC300_M0S0 1'b1
`else
	`define ATCBMC300_M0S0 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV1
	`define ATCBMC300_M0S1 1'b1
`else
	`define ATCBMC300_M0S1 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV2
	`define ATCBMC300_M0S2 1'b1
`else
	`define ATCBMC300_M0S2 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV3
	`define ATCBMC300_M0S3 1'b1
`else
	`define ATCBMC300_M0S3 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV4
	`define ATCBMC300_M0S4 1'b1
`else
	`define ATCBMC300_M0S4 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV5
	`define ATCBMC300_M0S5 1'b1
`else
	`define ATCBMC300_M0S5 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV6
	`define ATCBMC300_M0S6 1'b1
`else
	`define ATCBMC300_M0S6 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV7
	`define ATCBMC300_M0S7 1'b1
`else
	`define ATCBMC300_M0S7 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV8
	`define ATCBMC300_M0S8 1'b1
`else
	`define ATCBMC300_M0S8 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV9
	`define ATCBMC300_M0S9 1'b1
`else
	`define ATCBMC300_M0S9 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV10
	`define ATCBMC300_M0S10 1'b1
`else
	`define ATCBMC300_M0S10 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV11
	`define ATCBMC300_M0S11 1'b1
`else
	`define ATCBMC300_M0S11 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV12
	`define ATCBMC300_M0S12 1'b1
`else
	`define ATCBMC300_M0S12 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV13
	`define ATCBMC300_M0S13 1'b1
`else
	`define ATCBMC300_M0S13 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV14
	`define ATCBMC300_M0S14 1'b1
`else
	`define ATCBMC300_M0S14 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV15
	`define ATCBMC300_M0S15 1'b1
`else
	`define ATCBMC300_M0S15 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV16
	`define ATCBMC300_M0S16 1'b1
`else
	`define ATCBMC300_M0S16 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV17
	`define ATCBMC300_M0S17 1'b1
`else
	`define ATCBMC300_M0S17 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV18
	`define ATCBMC300_M0S18 1'b1
`else
	`define ATCBMC300_M0S18 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV19
	`define ATCBMC300_M0S19 1'b1
`else
	`define ATCBMC300_M0S19 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV20
	`define ATCBMC300_M0S20 1'b1
`else
	`define ATCBMC300_M0S20 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV21
	`define ATCBMC300_M0S21 1'b1
`else
	`define ATCBMC300_M0S21 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV22
	`define ATCBMC300_M0S22 1'b1
`else
	`define ATCBMC300_M0S22 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV23
	`define ATCBMC300_M0S23 1'b1
`else
	`define ATCBMC300_M0S23 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV24
	`define ATCBMC300_M0S24 1'b1
`else
	`define ATCBMC300_M0S24 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV25
	`define ATCBMC300_M0S25 1'b1
`else
	`define ATCBMC300_M0S25 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV26
	`define ATCBMC300_M0S26 1'b1
`else
	`define ATCBMC300_M0S26 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV27
	`define ATCBMC300_M0S27 1'b1
`else
	`define ATCBMC300_M0S27 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV28
	`define ATCBMC300_M0S28 1'b1
`else
	`define ATCBMC300_M0S28 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV29
	`define ATCBMC300_M0S29 1'b1
`else
	`define ATCBMC300_M0S29 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV30
	`define ATCBMC300_M0S30 1'b1
`else
	`define ATCBMC300_M0S30 1'b0
`endif
`ifdef ATCBMC300_MST0_SLV31
	`define ATCBMC300_M0S31 1'b1
`else
	`define ATCBMC300_M0S31 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV0
	`define ATCBMC300_M1S0 1'b1
`else
	`define ATCBMC300_M1S0 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV1
	`define ATCBMC300_M1S1 1'b1
`else
	`define ATCBMC300_M1S1 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV2
	`define ATCBMC300_M1S2 1'b1
`else
	`define ATCBMC300_M1S2 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV3
	`define ATCBMC300_M1S3 1'b1
`else
	`define ATCBMC300_M1S3 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV4
	`define ATCBMC300_M1S4 1'b1
`else
	`define ATCBMC300_M1S4 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV5
	`define ATCBMC300_M1S5 1'b1
`else
	`define ATCBMC300_M1S5 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV6
	`define ATCBMC300_M1S6 1'b1
`else
	`define ATCBMC300_M1S6 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV7
	`define ATCBMC300_M1S7 1'b1
`else
	`define ATCBMC300_M1S7 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV8
	`define ATCBMC300_M1S8 1'b1
`else
	`define ATCBMC300_M1S8 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV9
	`define ATCBMC300_M1S9 1'b1
`else
	`define ATCBMC300_M1S9 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV10
	`define ATCBMC300_M1S10 1'b1
`else
	`define ATCBMC300_M1S10 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV11
	`define ATCBMC300_M1S11 1'b1
`else
	`define ATCBMC300_M1S11 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV12
	`define ATCBMC300_M1S12 1'b1
`else
	`define ATCBMC300_M1S12 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV13
	`define ATCBMC300_M1S13 1'b1
`else
	`define ATCBMC300_M1S13 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV14
	`define ATCBMC300_M1S14 1'b1
`else
	`define ATCBMC300_M1S14 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV15
	`define ATCBMC300_M1S15 1'b1
`else
	`define ATCBMC300_M1S15 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV16
	`define ATCBMC300_M1S16 1'b1
`else
	`define ATCBMC300_M1S16 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV17
	`define ATCBMC300_M1S17 1'b1
`else
	`define ATCBMC300_M1S17 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV18
	`define ATCBMC300_M1S18 1'b1
`else
	`define ATCBMC300_M1S18 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV19
	`define ATCBMC300_M1S19 1'b1
`else
	`define ATCBMC300_M1S19 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV20
	`define ATCBMC300_M1S20 1'b1
`else
	`define ATCBMC300_M1S20 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV21
	`define ATCBMC300_M1S21 1'b1
`else
	`define ATCBMC300_M1S21 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV22
	`define ATCBMC300_M1S22 1'b1
`else
	`define ATCBMC300_M1S22 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV23
	`define ATCBMC300_M1S23 1'b1
`else
	`define ATCBMC300_M1S23 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV24
	`define ATCBMC300_M1S24 1'b1
`else
	`define ATCBMC300_M1S24 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV25
	`define ATCBMC300_M1S25 1'b1
`else
	`define ATCBMC300_M1S25 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV26
	`define ATCBMC300_M1S26 1'b1
`else
	`define ATCBMC300_M1S26 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV27
	`define ATCBMC300_M1S27 1'b1
`else
	`define ATCBMC300_M1S27 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV28
	`define ATCBMC300_M1S28 1'b1
`else
	`define ATCBMC300_M1S28 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV29
	`define ATCBMC300_M1S29 1'b1
`else
	`define ATCBMC300_M1S29 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV30
	`define ATCBMC300_M1S30 1'b1
`else
	`define ATCBMC300_M1S30 1'b0
`endif
`ifdef ATCBMC300_MST1_SLV31
	`define ATCBMC300_M1S31 1'b1
`else
	`define ATCBMC300_M1S31 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV0
	`define ATCBMC300_M2S0 1'b1
`else
	`define ATCBMC300_M2S0 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV1
	`define ATCBMC300_M2S1 1'b1
`else
	`define ATCBMC300_M2S1 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV2
	`define ATCBMC300_M2S2 1'b1
`else
	`define ATCBMC300_M2S2 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV3
	`define ATCBMC300_M2S3 1'b1
`else
	`define ATCBMC300_M2S3 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV4
	`define ATCBMC300_M2S4 1'b1
`else
	`define ATCBMC300_M2S4 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV5
	`define ATCBMC300_M2S5 1'b1
`else
	`define ATCBMC300_M2S5 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV6
	`define ATCBMC300_M2S6 1'b1
`else
	`define ATCBMC300_M2S6 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV7
	`define ATCBMC300_M2S7 1'b1
`else
	`define ATCBMC300_M2S7 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV8
	`define ATCBMC300_M2S8 1'b1
`else
	`define ATCBMC300_M2S8 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV9
	`define ATCBMC300_M2S9 1'b1
`else
	`define ATCBMC300_M2S9 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV10
	`define ATCBMC300_M2S10 1'b1
`else
	`define ATCBMC300_M2S10 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV11
	`define ATCBMC300_M2S11 1'b1
`else
	`define ATCBMC300_M2S11 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV12
	`define ATCBMC300_M2S12 1'b1
`else
	`define ATCBMC300_M2S12 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV13
	`define ATCBMC300_M2S13 1'b1
`else
	`define ATCBMC300_M2S13 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV14
	`define ATCBMC300_M2S14 1'b1
`else
	`define ATCBMC300_M2S14 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV15
	`define ATCBMC300_M2S15 1'b1
`else
	`define ATCBMC300_M2S15 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV16
	`define ATCBMC300_M2S16 1'b1
`else
	`define ATCBMC300_M2S16 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV17
	`define ATCBMC300_M2S17 1'b1
`else
	`define ATCBMC300_M2S17 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV18
	`define ATCBMC300_M2S18 1'b1
`else
	`define ATCBMC300_M2S18 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV19
	`define ATCBMC300_M2S19 1'b1
`else
	`define ATCBMC300_M2S19 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV20
	`define ATCBMC300_M2S20 1'b1
`else
	`define ATCBMC300_M2S20 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV21
	`define ATCBMC300_M2S21 1'b1
`else
	`define ATCBMC300_M2S21 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV22
	`define ATCBMC300_M2S22 1'b1
`else
	`define ATCBMC300_M2S22 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV23
	`define ATCBMC300_M2S23 1'b1
`else
	`define ATCBMC300_M2S23 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV24
	`define ATCBMC300_M2S24 1'b1
`else
	`define ATCBMC300_M2S24 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV25
	`define ATCBMC300_M2S25 1'b1
`else
	`define ATCBMC300_M2S25 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV26
	`define ATCBMC300_M2S26 1'b1
`else
	`define ATCBMC300_M2S26 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV27
	`define ATCBMC300_M2S27 1'b1
`else
	`define ATCBMC300_M2S27 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV28
	`define ATCBMC300_M2S28 1'b1
`else
	`define ATCBMC300_M2S28 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV29
	`define ATCBMC300_M2S29 1'b1
`else
	`define ATCBMC300_M2S29 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV30
	`define ATCBMC300_M2S30 1'b1
`else
	`define ATCBMC300_M2S30 1'b0
`endif
`ifdef ATCBMC300_MST2_SLV31
	`define ATCBMC300_M2S31 1'b1
`else
	`define ATCBMC300_M2S31 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV0
	`define ATCBMC300_M3S0 1'b1
`else
	`define ATCBMC300_M3S0 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV1
	`define ATCBMC300_M3S1 1'b1
`else
	`define ATCBMC300_M3S1 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV2
	`define ATCBMC300_M3S2 1'b1
`else
	`define ATCBMC300_M3S2 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV3
	`define ATCBMC300_M3S3 1'b1
`else
	`define ATCBMC300_M3S3 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV4
	`define ATCBMC300_M3S4 1'b1
`else
	`define ATCBMC300_M3S4 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV5
	`define ATCBMC300_M3S5 1'b1
`else
	`define ATCBMC300_M3S5 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV6
	`define ATCBMC300_M3S6 1'b1
`else
	`define ATCBMC300_M3S6 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV7
	`define ATCBMC300_M3S7 1'b1
`else
	`define ATCBMC300_M3S7 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV8
	`define ATCBMC300_M3S8 1'b1
`else
	`define ATCBMC300_M3S8 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV9
	`define ATCBMC300_M3S9 1'b1
`else
	`define ATCBMC300_M3S9 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV10
	`define ATCBMC300_M3S10 1'b1
`else
	`define ATCBMC300_M3S10 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV11
	`define ATCBMC300_M3S11 1'b1
`else
	`define ATCBMC300_M3S11 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV12
	`define ATCBMC300_M3S12 1'b1
`else
	`define ATCBMC300_M3S12 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV13
	`define ATCBMC300_M3S13 1'b1
`else
	`define ATCBMC300_M3S13 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV14
	`define ATCBMC300_M3S14 1'b1
`else
	`define ATCBMC300_M3S14 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV15
	`define ATCBMC300_M3S15 1'b1
`else
	`define ATCBMC300_M3S15 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV16
	`define ATCBMC300_M3S16 1'b1
`else
	`define ATCBMC300_M3S16 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV17
	`define ATCBMC300_M3S17 1'b1
`else
	`define ATCBMC300_M3S17 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV18
	`define ATCBMC300_M3S18 1'b1
`else
	`define ATCBMC300_M3S18 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV19
	`define ATCBMC300_M3S19 1'b1
`else
	`define ATCBMC300_M3S19 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV20
	`define ATCBMC300_M3S20 1'b1
`else
	`define ATCBMC300_M3S20 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV21
	`define ATCBMC300_M3S21 1'b1
`else
	`define ATCBMC300_M3S21 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV22
	`define ATCBMC300_M3S22 1'b1
`else
	`define ATCBMC300_M3S22 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV23
	`define ATCBMC300_M3S23 1'b1
`else
	`define ATCBMC300_M3S23 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV24
	`define ATCBMC300_M3S24 1'b1
`else
	`define ATCBMC300_M3S24 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV25
	`define ATCBMC300_M3S25 1'b1
`else
	`define ATCBMC300_M3S25 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV26
	`define ATCBMC300_M3S26 1'b1
`else
	`define ATCBMC300_M3S26 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV27
	`define ATCBMC300_M3S27 1'b1
`else
	`define ATCBMC300_M3S27 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV28
	`define ATCBMC300_M3S28 1'b1
`else
	`define ATCBMC300_M3S28 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV29
	`define ATCBMC300_M3S29 1'b1
`else
	`define ATCBMC300_M3S29 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV30
	`define ATCBMC300_M3S30 1'b1
`else
	`define ATCBMC300_M3S30 1'b0
`endif
`ifdef ATCBMC300_MST3_SLV31
	`define ATCBMC300_M3S31 1'b1
`else
	`define ATCBMC300_M3S31 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV0
	`define ATCBMC300_M4S0 1'b1
`else
	`define ATCBMC300_M4S0 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV1
	`define ATCBMC300_M4S1 1'b1
`else
	`define ATCBMC300_M4S1 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV2
	`define ATCBMC300_M4S2 1'b1
`else
	`define ATCBMC300_M4S2 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV3
	`define ATCBMC300_M4S3 1'b1
`else
	`define ATCBMC300_M4S3 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV4
	`define ATCBMC300_M4S4 1'b1
`else
	`define ATCBMC300_M4S4 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV5
	`define ATCBMC300_M4S5 1'b1
`else
	`define ATCBMC300_M4S5 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV6
	`define ATCBMC300_M4S6 1'b1
`else
	`define ATCBMC300_M4S6 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV7
	`define ATCBMC300_M4S7 1'b1
`else
	`define ATCBMC300_M4S7 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV8
	`define ATCBMC300_M4S8 1'b1
`else
	`define ATCBMC300_M4S8 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV9
	`define ATCBMC300_M4S9 1'b1
`else
	`define ATCBMC300_M4S9 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV10
	`define ATCBMC300_M4S10 1'b1
`else
	`define ATCBMC300_M4S10 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV11
	`define ATCBMC300_M4S11 1'b1
`else
	`define ATCBMC300_M4S11 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV12
	`define ATCBMC300_M4S12 1'b1
`else
	`define ATCBMC300_M4S12 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV13
	`define ATCBMC300_M4S13 1'b1
`else
	`define ATCBMC300_M4S13 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV14
	`define ATCBMC300_M4S14 1'b1
`else
	`define ATCBMC300_M4S14 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV15
	`define ATCBMC300_M4S15 1'b1
`else
	`define ATCBMC300_M4S15 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV16
	`define ATCBMC300_M4S16 1'b1
`else
	`define ATCBMC300_M4S16 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV17
	`define ATCBMC300_M4S17 1'b1
`else
	`define ATCBMC300_M4S17 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV18
	`define ATCBMC300_M4S18 1'b1
`else
	`define ATCBMC300_M4S18 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV19
	`define ATCBMC300_M4S19 1'b1
`else
	`define ATCBMC300_M4S19 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV20
	`define ATCBMC300_M4S20 1'b1
`else
	`define ATCBMC300_M4S20 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV21
	`define ATCBMC300_M4S21 1'b1
`else
	`define ATCBMC300_M4S21 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV22
	`define ATCBMC300_M4S22 1'b1
`else
	`define ATCBMC300_M4S22 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV23
	`define ATCBMC300_M4S23 1'b1
`else
	`define ATCBMC300_M4S23 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV24
	`define ATCBMC300_M4S24 1'b1
`else
	`define ATCBMC300_M4S24 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV25
	`define ATCBMC300_M4S25 1'b1
`else
	`define ATCBMC300_M4S25 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV26
	`define ATCBMC300_M4S26 1'b1
`else
	`define ATCBMC300_M4S26 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV27
	`define ATCBMC300_M4S27 1'b1
`else
	`define ATCBMC300_M4S27 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV28
	`define ATCBMC300_M4S28 1'b1
`else
	`define ATCBMC300_M4S28 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV29
	`define ATCBMC300_M4S29 1'b1
`else
	`define ATCBMC300_M4S29 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV30
	`define ATCBMC300_M4S30 1'b1
`else
	`define ATCBMC300_M4S30 1'b0
`endif
`ifdef ATCBMC300_MST4_SLV31
	`define ATCBMC300_M4S31 1'b1
`else
	`define ATCBMC300_M4S31 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV0
	`define ATCBMC300_M5S0 1'b1
`else
	`define ATCBMC300_M5S0 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV1
	`define ATCBMC300_M5S1 1'b1
`else
	`define ATCBMC300_M5S1 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV2
	`define ATCBMC300_M5S2 1'b1
`else
	`define ATCBMC300_M5S2 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV3
	`define ATCBMC300_M5S3 1'b1
`else
	`define ATCBMC300_M5S3 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV4
	`define ATCBMC300_M5S4 1'b1
`else
	`define ATCBMC300_M5S4 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV5
	`define ATCBMC300_M5S5 1'b1
`else
	`define ATCBMC300_M5S5 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV6
	`define ATCBMC300_M5S6 1'b1
`else
	`define ATCBMC300_M5S6 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV7
	`define ATCBMC300_M5S7 1'b1
`else
	`define ATCBMC300_M5S7 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV8
	`define ATCBMC300_M5S8 1'b1
`else
	`define ATCBMC300_M5S8 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV9
	`define ATCBMC300_M5S9 1'b1
`else
	`define ATCBMC300_M5S9 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV10
	`define ATCBMC300_M5S10 1'b1
`else
	`define ATCBMC300_M5S10 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV11
	`define ATCBMC300_M5S11 1'b1
`else
	`define ATCBMC300_M5S11 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV12
	`define ATCBMC300_M5S12 1'b1
`else
	`define ATCBMC300_M5S12 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV13
	`define ATCBMC300_M5S13 1'b1
`else
	`define ATCBMC300_M5S13 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV14
	`define ATCBMC300_M5S14 1'b1
`else
	`define ATCBMC300_M5S14 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV15
	`define ATCBMC300_M5S15 1'b1
`else
	`define ATCBMC300_M5S15 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV16
	`define ATCBMC300_M5S16 1'b1
`else
	`define ATCBMC300_M5S16 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV17
	`define ATCBMC300_M5S17 1'b1
`else
	`define ATCBMC300_M5S17 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV18
	`define ATCBMC300_M5S18 1'b1
`else
	`define ATCBMC300_M5S18 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV19
	`define ATCBMC300_M5S19 1'b1
`else
	`define ATCBMC300_M5S19 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV20
	`define ATCBMC300_M5S20 1'b1
`else
	`define ATCBMC300_M5S20 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV21
	`define ATCBMC300_M5S21 1'b1
`else
	`define ATCBMC300_M5S21 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV22
	`define ATCBMC300_M5S22 1'b1
`else
	`define ATCBMC300_M5S22 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV23
	`define ATCBMC300_M5S23 1'b1
`else
	`define ATCBMC300_M5S23 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV24
	`define ATCBMC300_M5S24 1'b1
`else
	`define ATCBMC300_M5S24 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV25
	`define ATCBMC300_M5S25 1'b1
`else
	`define ATCBMC300_M5S25 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV26
	`define ATCBMC300_M5S26 1'b1
`else
	`define ATCBMC300_M5S26 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV27
	`define ATCBMC300_M5S27 1'b1
`else
	`define ATCBMC300_M5S27 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV28
	`define ATCBMC300_M5S28 1'b1
`else
	`define ATCBMC300_M5S28 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV29
	`define ATCBMC300_M5S29 1'b1
`else
	`define ATCBMC300_M5S29 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV30
	`define ATCBMC300_M5S30 1'b1
`else
	`define ATCBMC300_M5S30 1'b0
`endif
`ifdef ATCBMC300_MST5_SLV31
	`define ATCBMC300_M5S31 1'b1
`else
	`define ATCBMC300_M5S31 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV0
	`define ATCBMC300_M6S0 1'b1
`else
	`define ATCBMC300_M6S0 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV1
	`define ATCBMC300_M6S1 1'b1
`else
	`define ATCBMC300_M6S1 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV2
	`define ATCBMC300_M6S2 1'b1
`else
	`define ATCBMC300_M6S2 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV3
	`define ATCBMC300_M6S3 1'b1
`else
	`define ATCBMC300_M6S3 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV4
	`define ATCBMC300_M6S4 1'b1
`else
	`define ATCBMC300_M6S4 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV5
	`define ATCBMC300_M6S5 1'b1
`else
	`define ATCBMC300_M6S5 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV6
	`define ATCBMC300_M6S6 1'b1
`else
	`define ATCBMC300_M6S6 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV7
	`define ATCBMC300_M6S7 1'b1
`else
	`define ATCBMC300_M6S7 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV8
	`define ATCBMC300_M6S8 1'b1
`else
	`define ATCBMC300_M6S8 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV9
	`define ATCBMC300_M6S9 1'b1
`else
	`define ATCBMC300_M6S9 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV10
	`define ATCBMC300_M6S10 1'b1
`else
	`define ATCBMC300_M6S10 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV11
	`define ATCBMC300_M6S11 1'b1
`else
	`define ATCBMC300_M6S11 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV12
	`define ATCBMC300_M6S12 1'b1
`else
	`define ATCBMC300_M6S12 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV13
	`define ATCBMC300_M6S13 1'b1
`else
	`define ATCBMC300_M6S13 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV14
	`define ATCBMC300_M6S14 1'b1
`else
	`define ATCBMC300_M6S14 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV15
	`define ATCBMC300_M6S15 1'b1
`else
	`define ATCBMC300_M6S15 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV16
	`define ATCBMC300_M6S16 1'b1
`else
	`define ATCBMC300_M6S16 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV17
	`define ATCBMC300_M6S17 1'b1
`else
	`define ATCBMC300_M6S17 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV18
	`define ATCBMC300_M6S18 1'b1
`else
	`define ATCBMC300_M6S18 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV19
	`define ATCBMC300_M6S19 1'b1
`else
	`define ATCBMC300_M6S19 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV20
	`define ATCBMC300_M6S20 1'b1
`else
	`define ATCBMC300_M6S20 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV21
	`define ATCBMC300_M6S21 1'b1
`else
	`define ATCBMC300_M6S21 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV22
	`define ATCBMC300_M6S22 1'b1
`else
	`define ATCBMC300_M6S22 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV23
	`define ATCBMC300_M6S23 1'b1
`else
	`define ATCBMC300_M6S23 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV24
	`define ATCBMC300_M6S24 1'b1
`else
	`define ATCBMC300_M6S24 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV25
	`define ATCBMC300_M6S25 1'b1
`else
	`define ATCBMC300_M6S25 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV26
	`define ATCBMC300_M6S26 1'b1
`else
	`define ATCBMC300_M6S26 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV27
	`define ATCBMC300_M6S27 1'b1
`else
	`define ATCBMC300_M6S27 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV28
	`define ATCBMC300_M6S28 1'b1
`else
	`define ATCBMC300_M6S28 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV29
	`define ATCBMC300_M6S29 1'b1
`else
	`define ATCBMC300_M6S29 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV30
	`define ATCBMC300_M6S30 1'b1
`else
	`define ATCBMC300_M6S30 1'b0
`endif
`ifdef ATCBMC300_MST6_SLV31
	`define ATCBMC300_M6S31 1'b1
`else
	`define ATCBMC300_M6S31 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV0
	`define ATCBMC300_M7S0 1'b1
`else
	`define ATCBMC300_M7S0 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV1
	`define ATCBMC300_M7S1 1'b1
`else
	`define ATCBMC300_M7S1 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV2
	`define ATCBMC300_M7S2 1'b1
`else
	`define ATCBMC300_M7S2 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV3
	`define ATCBMC300_M7S3 1'b1
`else
	`define ATCBMC300_M7S3 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV4
	`define ATCBMC300_M7S4 1'b1
`else
	`define ATCBMC300_M7S4 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV5
	`define ATCBMC300_M7S5 1'b1
`else
	`define ATCBMC300_M7S5 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV6
	`define ATCBMC300_M7S6 1'b1
`else
	`define ATCBMC300_M7S6 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV7
	`define ATCBMC300_M7S7 1'b1
`else
	`define ATCBMC300_M7S7 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV8
	`define ATCBMC300_M7S8 1'b1
`else
	`define ATCBMC300_M7S8 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV9
	`define ATCBMC300_M7S9 1'b1
`else
	`define ATCBMC300_M7S9 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV10
	`define ATCBMC300_M7S10 1'b1
`else
	`define ATCBMC300_M7S10 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV11
	`define ATCBMC300_M7S11 1'b1
`else
	`define ATCBMC300_M7S11 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV12
	`define ATCBMC300_M7S12 1'b1
`else
	`define ATCBMC300_M7S12 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV13
	`define ATCBMC300_M7S13 1'b1
`else
	`define ATCBMC300_M7S13 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV14
	`define ATCBMC300_M7S14 1'b1
`else
	`define ATCBMC300_M7S14 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV15
	`define ATCBMC300_M7S15 1'b1
`else
	`define ATCBMC300_M7S15 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV16
	`define ATCBMC300_M7S16 1'b1
`else
	`define ATCBMC300_M7S16 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV17
	`define ATCBMC300_M7S17 1'b1
`else
	`define ATCBMC300_M7S17 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV18
	`define ATCBMC300_M7S18 1'b1
`else
	`define ATCBMC300_M7S18 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV19
	`define ATCBMC300_M7S19 1'b1
`else
	`define ATCBMC300_M7S19 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV20
	`define ATCBMC300_M7S20 1'b1
`else
	`define ATCBMC300_M7S20 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV21
	`define ATCBMC300_M7S21 1'b1
`else
	`define ATCBMC300_M7S21 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV22
	`define ATCBMC300_M7S22 1'b1
`else
	`define ATCBMC300_M7S22 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV23
	`define ATCBMC300_M7S23 1'b1
`else
	`define ATCBMC300_M7S23 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV24
	`define ATCBMC300_M7S24 1'b1
`else
	`define ATCBMC300_M7S24 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV25
	`define ATCBMC300_M7S25 1'b1
`else
	`define ATCBMC300_M7S25 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV26
	`define ATCBMC300_M7S26 1'b1
`else
	`define ATCBMC300_M7S26 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV27
	`define ATCBMC300_M7S27 1'b1
`else
	`define ATCBMC300_M7S27 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV28
	`define ATCBMC300_M7S28 1'b1
`else
	`define ATCBMC300_M7S28 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV29
	`define ATCBMC300_M7S29 1'b1
`else
	`define ATCBMC300_M7S29 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV30
	`define ATCBMC300_M7S30 1'b1
`else
	`define ATCBMC300_M7S30 1'b0
`endif
`ifdef ATCBMC300_MST7_SLV31
	`define ATCBMC300_M7S31 1'b1
`else
	`define ATCBMC300_M7S31 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV0
	`define ATCBMC300_M8S0 1'b1
`else
	`define ATCBMC300_M8S0 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV1
	`define ATCBMC300_M8S1 1'b1
`else
	`define ATCBMC300_M8S1 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV2
	`define ATCBMC300_M8S2 1'b1
`else
	`define ATCBMC300_M8S2 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV3
	`define ATCBMC300_M8S3 1'b1
`else
	`define ATCBMC300_M8S3 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV4
	`define ATCBMC300_M8S4 1'b1
`else
	`define ATCBMC300_M8S4 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV5
	`define ATCBMC300_M8S5 1'b1
`else
	`define ATCBMC300_M8S5 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV6
	`define ATCBMC300_M8S6 1'b1
`else
	`define ATCBMC300_M8S6 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV7
	`define ATCBMC300_M8S7 1'b1
`else
	`define ATCBMC300_M8S7 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV8
	`define ATCBMC300_M8S8 1'b1
`else
	`define ATCBMC300_M8S8 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV9
	`define ATCBMC300_M8S9 1'b1
`else
	`define ATCBMC300_M8S9 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV10
	`define ATCBMC300_M8S10 1'b1
`else
	`define ATCBMC300_M8S10 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV11
	`define ATCBMC300_M8S11 1'b1
`else
	`define ATCBMC300_M8S11 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV12
	`define ATCBMC300_M8S12 1'b1
`else
	`define ATCBMC300_M8S12 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV13
	`define ATCBMC300_M8S13 1'b1
`else
	`define ATCBMC300_M8S13 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV14
	`define ATCBMC300_M8S14 1'b1
`else
	`define ATCBMC300_M8S14 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV15
	`define ATCBMC300_M8S15 1'b1
`else
	`define ATCBMC300_M8S15 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV16
	`define ATCBMC300_M8S16 1'b1
`else
	`define ATCBMC300_M8S16 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV17
	`define ATCBMC300_M8S17 1'b1
`else
	`define ATCBMC300_M8S17 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV18
	`define ATCBMC300_M8S18 1'b1
`else
	`define ATCBMC300_M8S18 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV19
	`define ATCBMC300_M8S19 1'b1
`else
	`define ATCBMC300_M8S19 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV20
	`define ATCBMC300_M8S20 1'b1
`else
	`define ATCBMC300_M8S20 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV21
	`define ATCBMC300_M8S21 1'b1
`else
	`define ATCBMC300_M8S21 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV22
	`define ATCBMC300_M8S22 1'b1
`else
	`define ATCBMC300_M8S22 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV23
	`define ATCBMC300_M8S23 1'b1
`else
	`define ATCBMC300_M8S23 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV24
	`define ATCBMC300_M8S24 1'b1
`else
	`define ATCBMC300_M8S24 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV25
	`define ATCBMC300_M8S25 1'b1
`else
	`define ATCBMC300_M8S25 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV26
	`define ATCBMC300_M8S26 1'b1
`else
	`define ATCBMC300_M8S26 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV27
	`define ATCBMC300_M8S27 1'b1
`else
	`define ATCBMC300_M8S27 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV28
	`define ATCBMC300_M8S28 1'b1
`else
	`define ATCBMC300_M8S28 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV29
	`define ATCBMC300_M8S29 1'b1
`else
	`define ATCBMC300_M8S29 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV30
	`define ATCBMC300_M8S30 1'b1
`else
	`define ATCBMC300_M8S30 1'b0
`endif
`ifdef ATCBMC300_MST8_SLV31
	`define ATCBMC300_M8S31 1'b1
`else
	`define ATCBMC300_M8S31 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV0
	`define ATCBMC300_M9S0 1'b1
`else
	`define ATCBMC300_M9S0 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV1
	`define ATCBMC300_M9S1 1'b1
`else
	`define ATCBMC300_M9S1 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV2
	`define ATCBMC300_M9S2 1'b1
`else
	`define ATCBMC300_M9S2 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV3
	`define ATCBMC300_M9S3 1'b1
`else
	`define ATCBMC300_M9S3 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV4
	`define ATCBMC300_M9S4 1'b1
`else
	`define ATCBMC300_M9S4 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV5
	`define ATCBMC300_M9S5 1'b1
`else
	`define ATCBMC300_M9S5 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV6
	`define ATCBMC300_M9S6 1'b1
`else
	`define ATCBMC300_M9S6 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV7
	`define ATCBMC300_M9S7 1'b1
`else
	`define ATCBMC300_M9S7 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV8
	`define ATCBMC300_M9S8 1'b1
`else
	`define ATCBMC300_M9S8 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV9
	`define ATCBMC300_M9S9 1'b1
`else
	`define ATCBMC300_M9S9 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV10
	`define ATCBMC300_M9S10 1'b1
`else
	`define ATCBMC300_M9S10 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV11
	`define ATCBMC300_M9S11 1'b1
`else
	`define ATCBMC300_M9S11 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV12
	`define ATCBMC300_M9S12 1'b1
`else
	`define ATCBMC300_M9S12 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV13
	`define ATCBMC300_M9S13 1'b1
`else
	`define ATCBMC300_M9S13 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV14
	`define ATCBMC300_M9S14 1'b1
`else
	`define ATCBMC300_M9S14 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV15
	`define ATCBMC300_M9S15 1'b1
`else
	`define ATCBMC300_M9S15 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV16
	`define ATCBMC300_M9S16 1'b1
`else
	`define ATCBMC300_M9S16 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV17
	`define ATCBMC300_M9S17 1'b1
`else
	`define ATCBMC300_M9S17 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV18
	`define ATCBMC300_M9S18 1'b1
`else
	`define ATCBMC300_M9S18 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV19
	`define ATCBMC300_M9S19 1'b1
`else
	`define ATCBMC300_M9S19 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV20
	`define ATCBMC300_M9S20 1'b1
`else
	`define ATCBMC300_M9S20 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV21
	`define ATCBMC300_M9S21 1'b1
`else
	`define ATCBMC300_M9S21 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV22
	`define ATCBMC300_M9S22 1'b1
`else
	`define ATCBMC300_M9S22 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV23
	`define ATCBMC300_M9S23 1'b1
`else
	`define ATCBMC300_M9S23 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV24
	`define ATCBMC300_M9S24 1'b1
`else
	`define ATCBMC300_M9S24 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV25
	`define ATCBMC300_M9S25 1'b1
`else
	`define ATCBMC300_M9S25 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV26
	`define ATCBMC300_M9S26 1'b1
`else
	`define ATCBMC300_M9S26 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV27
	`define ATCBMC300_M9S27 1'b1
`else
	`define ATCBMC300_M9S27 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV28
	`define ATCBMC300_M9S28 1'b1
`else
	`define ATCBMC300_M9S28 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV29
	`define ATCBMC300_M9S29 1'b1
`else
	`define ATCBMC300_M9S29 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV30
	`define ATCBMC300_M9S30 1'b1
`else
	`define ATCBMC300_M9S30 1'b0
`endif
`ifdef ATCBMC300_MST9_SLV31
	`define ATCBMC300_M9S31 1'b1
`else
	`define ATCBMC300_M9S31 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV0
	`define ATCBMC300_M10S0 1'b1
`else
	`define ATCBMC300_M10S0 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV1
	`define ATCBMC300_M10S1 1'b1
`else
	`define ATCBMC300_M10S1 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV2
	`define ATCBMC300_M10S2 1'b1
`else
	`define ATCBMC300_M10S2 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV3
	`define ATCBMC300_M10S3 1'b1
`else
	`define ATCBMC300_M10S3 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV4
	`define ATCBMC300_M10S4 1'b1
`else
	`define ATCBMC300_M10S4 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV5
	`define ATCBMC300_M10S5 1'b1
`else
	`define ATCBMC300_M10S5 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV6
	`define ATCBMC300_M10S6 1'b1
`else
	`define ATCBMC300_M10S6 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV7
	`define ATCBMC300_M10S7 1'b1
`else
	`define ATCBMC300_M10S7 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV8
	`define ATCBMC300_M10S8 1'b1
`else
	`define ATCBMC300_M10S8 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV9
	`define ATCBMC300_M10S9 1'b1
`else
	`define ATCBMC300_M10S9 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV10
	`define ATCBMC300_M10S10 1'b1
`else
	`define ATCBMC300_M10S10 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV11
	`define ATCBMC300_M10S11 1'b1
`else
	`define ATCBMC300_M10S11 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV12
	`define ATCBMC300_M10S12 1'b1
`else
	`define ATCBMC300_M10S12 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV13
	`define ATCBMC300_M10S13 1'b1
`else
	`define ATCBMC300_M10S13 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV14
	`define ATCBMC300_M10S14 1'b1
`else
	`define ATCBMC300_M10S14 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV15
	`define ATCBMC300_M10S15 1'b1
`else
	`define ATCBMC300_M10S15 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV16
	`define ATCBMC300_M10S16 1'b1
`else
	`define ATCBMC300_M10S16 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV17
	`define ATCBMC300_M10S17 1'b1
`else
	`define ATCBMC300_M10S17 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV18
	`define ATCBMC300_M10S18 1'b1
`else
	`define ATCBMC300_M10S18 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV19
	`define ATCBMC300_M10S19 1'b1
`else
	`define ATCBMC300_M10S19 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV20
	`define ATCBMC300_M10S20 1'b1
`else
	`define ATCBMC300_M10S20 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV21
	`define ATCBMC300_M10S21 1'b1
`else
	`define ATCBMC300_M10S21 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV22
	`define ATCBMC300_M10S22 1'b1
`else
	`define ATCBMC300_M10S22 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV23
	`define ATCBMC300_M10S23 1'b1
`else
	`define ATCBMC300_M10S23 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV24
	`define ATCBMC300_M10S24 1'b1
`else
	`define ATCBMC300_M10S24 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV25
	`define ATCBMC300_M10S25 1'b1
`else
	`define ATCBMC300_M10S25 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV26
	`define ATCBMC300_M10S26 1'b1
`else
	`define ATCBMC300_M10S26 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV27
	`define ATCBMC300_M10S27 1'b1
`else
	`define ATCBMC300_M10S27 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV28
	`define ATCBMC300_M10S28 1'b1
`else
	`define ATCBMC300_M10S28 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV29
	`define ATCBMC300_M10S29 1'b1
`else
	`define ATCBMC300_M10S29 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV30
	`define ATCBMC300_M10S30 1'b1
`else
	`define ATCBMC300_M10S30 1'b0
`endif
`ifdef ATCBMC300_MST10_SLV31
	`define ATCBMC300_M10S31 1'b1
`else
	`define ATCBMC300_M10S31 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV0
	`define ATCBMC300_M11S0 1'b1
`else
	`define ATCBMC300_M11S0 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV1
	`define ATCBMC300_M11S1 1'b1
`else
	`define ATCBMC300_M11S1 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV2
	`define ATCBMC300_M11S2 1'b1
`else
	`define ATCBMC300_M11S2 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV3
	`define ATCBMC300_M11S3 1'b1
`else
	`define ATCBMC300_M11S3 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV4
	`define ATCBMC300_M11S4 1'b1
`else
	`define ATCBMC300_M11S4 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV5
	`define ATCBMC300_M11S5 1'b1
`else
	`define ATCBMC300_M11S5 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV6
	`define ATCBMC300_M11S6 1'b1
`else
	`define ATCBMC300_M11S6 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV7
	`define ATCBMC300_M11S7 1'b1
`else
	`define ATCBMC300_M11S7 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV8
	`define ATCBMC300_M11S8 1'b1
`else
	`define ATCBMC300_M11S8 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV9
	`define ATCBMC300_M11S9 1'b1
`else
	`define ATCBMC300_M11S9 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV10
	`define ATCBMC300_M11S10 1'b1
`else
	`define ATCBMC300_M11S10 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV11
	`define ATCBMC300_M11S11 1'b1
`else
	`define ATCBMC300_M11S11 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV12
	`define ATCBMC300_M11S12 1'b1
`else
	`define ATCBMC300_M11S12 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV13
	`define ATCBMC300_M11S13 1'b1
`else
	`define ATCBMC300_M11S13 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV14
	`define ATCBMC300_M11S14 1'b1
`else
	`define ATCBMC300_M11S14 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV15
	`define ATCBMC300_M11S15 1'b1
`else
	`define ATCBMC300_M11S15 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV16
	`define ATCBMC300_M11S16 1'b1
`else
	`define ATCBMC300_M11S16 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV17
	`define ATCBMC300_M11S17 1'b1
`else
	`define ATCBMC300_M11S17 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV18
	`define ATCBMC300_M11S18 1'b1
`else
	`define ATCBMC300_M11S18 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV19
	`define ATCBMC300_M11S19 1'b1
`else
	`define ATCBMC300_M11S19 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV20
	`define ATCBMC300_M11S20 1'b1
`else
	`define ATCBMC300_M11S20 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV21
	`define ATCBMC300_M11S21 1'b1
`else
	`define ATCBMC300_M11S21 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV22
	`define ATCBMC300_M11S22 1'b1
`else
	`define ATCBMC300_M11S22 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV23
	`define ATCBMC300_M11S23 1'b1
`else
	`define ATCBMC300_M11S23 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV24
	`define ATCBMC300_M11S24 1'b1
`else
	`define ATCBMC300_M11S24 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV25
	`define ATCBMC300_M11S25 1'b1
`else
	`define ATCBMC300_M11S25 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV26
	`define ATCBMC300_M11S26 1'b1
`else
	`define ATCBMC300_M11S26 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV27
	`define ATCBMC300_M11S27 1'b1
`else
	`define ATCBMC300_M11S27 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV28
	`define ATCBMC300_M11S28 1'b1
`else
	`define ATCBMC300_M11S28 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV29
	`define ATCBMC300_M11S29 1'b1
`else
	`define ATCBMC300_M11S29 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV30
	`define ATCBMC300_M11S30 1'b1
`else
	`define ATCBMC300_M11S30 1'b0
`endif
`ifdef ATCBMC300_MST11_SLV31
	`define ATCBMC300_M11S31 1'b1
`else
	`define ATCBMC300_M11S31 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV0
	`define ATCBMC300_M12S0 1'b1
`else
	`define ATCBMC300_M12S0 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV1
	`define ATCBMC300_M12S1 1'b1
`else
	`define ATCBMC300_M12S1 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV2
	`define ATCBMC300_M12S2 1'b1
`else
	`define ATCBMC300_M12S2 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV3
	`define ATCBMC300_M12S3 1'b1
`else
	`define ATCBMC300_M12S3 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV4
	`define ATCBMC300_M12S4 1'b1
`else
	`define ATCBMC300_M12S4 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV5
	`define ATCBMC300_M12S5 1'b1
`else
	`define ATCBMC300_M12S5 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV6
	`define ATCBMC300_M12S6 1'b1
`else
	`define ATCBMC300_M12S6 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV7
	`define ATCBMC300_M12S7 1'b1
`else
	`define ATCBMC300_M12S7 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV8
	`define ATCBMC300_M12S8 1'b1
`else
	`define ATCBMC300_M12S8 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV9
	`define ATCBMC300_M12S9 1'b1
`else
	`define ATCBMC300_M12S9 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV10
	`define ATCBMC300_M12S10 1'b1
`else
	`define ATCBMC300_M12S10 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV11
	`define ATCBMC300_M12S11 1'b1
`else
	`define ATCBMC300_M12S11 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV12
	`define ATCBMC300_M12S12 1'b1
`else
	`define ATCBMC300_M12S12 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV13
	`define ATCBMC300_M12S13 1'b1
`else
	`define ATCBMC300_M12S13 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV14
	`define ATCBMC300_M12S14 1'b1
`else
	`define ATCBMC300_M12S14 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV15
	`define ATCBMC300_M12S15 1'b1
`else
	`define ATCBMC300_M12S15 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV16
	`define ATCBMC300_M12S16 1'b1
`else
	`define ATCBMC300_M12S16 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV17
	`define ATCBMC300_M12S17 1'b1
`else
	`define ATCBMC300_M12S17 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV18
	`define ATCBMC300_M12S18 1'b1
`else
	`define ATCBMC300_M12S18 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV19
	`define ATCBMC300_M12S19 1'b1
`else
	`define ATCBMC300_M12S19 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV20
	`define ATCBMC300_M12S20 1'b1
`else
	`define ATCBMC300_M12S20 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV21
	`define ATCBMC300_M12S21 1'b1
`else
	`define ATCBMC300_M12S21 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV22
	`define ATCBMC300_M12S22 1'b1
`else
	`define ATCBMC300_M12S22 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV23
	`define ATCBMC300_M12S23 1'b1
`else
	`define ATCBMC300_M12S23 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV24
	`define ATCBMC300_M12S24 1'b1
`else
	`define ATCBMC300_M12S24 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV25
	`define ATCBMC300_M12S25 1'b1
`else
	`define ATCBMC300_M12S25 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV26
	`define ATCBMC300_M12S26 1'b1
`else
	`define ATCBMC300_M12S26 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV27
	`define ATCBMC300_M12S27 1'b1
`else
	`define ATCBMC300_M12S27 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV28
	`define ATCBMC300_M12S28 1'b1
`else
	`define ATCBMC300_M12S28 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV29
	`define ATCBMC300_M12S29 1'b1
`else
	`define ATCBMC300_M12S29 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV30
	`define ATCBMC300_M12S30 1'b1
`else
	`define ATCBMC300_M12S30 1'b0
`endif
`ifdef ATCBMC300_MST12_SLV31
	`define ATCBMC300_M12S31 1'b1
`else
	`define ATCBMC300_M12S31 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV0
	`define ATCBMC300_M13S0 1'b1
`else
	`define ATCBMC300_M13S0 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV1
	`define ATCBMC300_M13S1 1'b1
`else
	`define ATCBMC300_M13S1 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV2
	`define ATCBMC300_M13S2 1'b1
`else
	`define ATCBMC300_M13S2 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV3
	`define ATCBMC300_M13S3 1'b1
`else
	`define ATCBMC300_M13S3 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV4
	`define ATCBMC300_M13S4 1'b1
`else
	`define ATCBMC300_M13S4 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV5
	`define ATCBMC300_M13S5 1'b1
`else
	`define ATCBMC300_M13S5 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV6
	`define ATCBMC300_M13S6 1'b1
`else
	`define ATCBMC300_M13S6 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV7
	`define ATCBMC300_M13S7 1'b1
`else
	`define ATCBMC300_M13S7 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV8
	`define ATCBMC300_M13S8 1'b1
`else
	`define ATCBMC300_M13S8 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV9
	`define ATCBMC300_M13S9 1'b1
`else
	`define ATCBMC300_M13S9 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV10
	`define ATCBMC300_M13S10 1'b1
`else
	`define ATCBMC300_M13S10 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV11
	`define ATCBMC300_M13S11 1'b1
`else
	`define ATCBMC300_M13S11 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV12
	`define ATCBMC300_M13S12 1'b1
`else
	`define ATCBMC300_M13S12 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV13
	`define ATCBMC300_M13S13 1'b1
`else
	`define ATCBMC300_M13S13 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV14
	`define ATCBMC300_M13S14 1'b1
`else
	`define ATCBMC300_M13S14 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV15
	`define ATCBMC300_M13S15 1'b1
`else
	`define ATCBMC300_M13S15 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV16
	`define ATCBMC300_M13S16 1'b1
`else
	`define ATCBMC300_M13S16 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV17
	`define ATCBMC300_M13S17 1'b1
`else
	`define ATCBMC300_M13S17 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV18
	`define ATCBMC300_M13S18 1'b1
`else
	`define ATCBMC300_M13S18 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV19
	`define ATCBMC300_M13S19 1'b1
`else
	`define ATCBMC300_M13S19 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV20
	`define ATCBMC300_M13S20 1'b1
`else
	`define ATCBMC300_M13S20 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV21
	`define ATCBMC300_M13S21 1'b1
`else
	`define ATCBMC300_M13S21 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV22
	`define ATCBMC300_M13S22 1'b1
`else
	`define ATCBMC300_M13S22 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV23
	`define ATCBMC300_M13S23 1'b1
`else
	`define ATCBMC300_M13S23 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV24
	`define ATCBMC300_M13S24 1'b1
`else
	`define ATCBMC300_M13S24 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV25
	`define ATCBMC300_M13S25 1'b1
`else
	`define ATCBMC300_M13S25 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV26
	`define ATCBMC300_M13S26 1'b1
`else
	`define ATCBMC300_M13S26 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV27
	`define ATCBMC300_M13S27 1'b1
`else
	`define ATCBMC300_M13S27 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV28
	`define ATCBMC300_M13S28 1'b1
`else
	`define ATCBMC300_M13S28 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV29
	`define ATCBMC300_M13S29 1'b1
`else
	`define ATCBMC300_M13S29 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV30
	`define ATCBMC300_M13S30 1'b1
`else
	`define ATCBMC300_M13S30 1'b0
`endif
`ifdef ATCBMC300_MST13_SLV31
	`define ATCBMC300_M13S31 1'b1
`else
	`define ATCBMC300_M13S31 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV0
	`define ATCBMC300_M14S0 1'b1
`else
	`define ATCBMC300_M14S0 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV1
	`define ATCBMC300_M14S1 1'b1
`else
	`define ATCBMC300_M14S1 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV2
	`define ATCBMC300_M14S2 1'b1
`else
	`define ATCBMC300_M14S2 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV3
	`define ATCBMC300_M14S3 1'b1
`else
	`define ATCBMC300_M14S3 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV4
	`define ATCBMC300_M14S4 1'b1
`else
	`define ATCBMC300_M14S4 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV5
	`define ATCBMC300_M14S5 1'b1
`else
	`define ATCBMC300_M14S5 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV6
	`define ATCBMC300_M14S6 1'b1
`else
	`define ATCBMC300_M14S6 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV7
	`define ATCBMC300_M14S7 1'b1
`else
	`define ATCBMC300_M14S7 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV8
	`define ATCBMC300_M14S8 1'b1
`else
	`define ATCBMC300_M14S8 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV9
	`define ATCBMC300_M14S9 1'b1
`else
	`define ATCBMC300_M14S9 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV10
	`define ATCBMC300_M14S10 1'b1
`else
	`define ATCBMC300_M14S10 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV11
	`define ATCBMC300_M14S11 1'b1
`else
	`define ATCBMC300_M14S11 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV12
	`define ATCBMC300_M14S12 1'b1
`else
	`define ATCBMC300_M14S12 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV13
	`define ATCBMC300_M14S13 1'b1
`else
	`define ATCBMC300_M14S13 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV14
	`define ATCBMC300_M14S14 1'b1
`else
	`define ATCBMC300_M14S14 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV15
	`define ATCBMC300_M14S15 1'b1
`else
	`define ATCBMC300_M14S15 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV16
	`define ATCBMC300_M14S16 1'b1
`else
	`define ATCBMC300_M14S16 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV17
	`define ATCBMC300_M14S17 1'b1
`else
	`define ATCBMC300_M14S17 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV18
	`define ATCBMC300_M14S18 1'b1
`else
	`define ATCBMC300_M14S18 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV19
	`define ATCBMC300_M14S19 1'b1
`else
	`define ATCBMC300_M14S19 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV20
	`define ATCBMC300_M14S20 1'b1
`else
	`define ATCBMC300_M14S20 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV21
	`define ATCBMC300_M14S21 1'b1
`else
	`define ATCBMC300_M14S21 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV22
	`define ATCBMC300_M14S22 1'b1
`else
	`define ATCBMC300_M14S22 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV23
	`define ATCBMC300_M14S23 1'b1
`else
	`define ATCBMC300_M14S23 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV24
	`define ATCBMC300_M14S24 1'b1
`else
	`define ATCBMC300_M14S24 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV25
	`define ATCBMC300_M14S25 1'b1
`else
	`define ATCBMC300_M14S25 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV26
	`define ATCBMC300_M14S26 1'b1
`else
	`define ATCBMC300_M14S26 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV27
	`define ATCBMC300_M14S27 1'b1
`else
	`define ATCBMC300_M14S27 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV28
	`define ATCBMC300_M14S28 1'b1
`else
	`define ATCBMC300_M14S28 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV29
	`define ATCBMC300_M14S29 1'b1
`else
	`define ATCBMC300_M14S29 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV30
	`define ATCBMC300_M14S30 1'b1
`else
	`define ATCBMC300_M14S30 1'b0
`endif
`ifdef ATCBMC300_MST14_SLV31
	`define ATCBMC300_M14S31 1'b1
`else
	`define ATCBMC300_M14S31 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV0
	`define ATCBMC300_M15S0 1'b1
`else
	`define ATCBMC300_M15S0 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV1
	`define ATCBMC300_M15S1 1'b1
`else
	`define ATCBMC300_M15S1 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV2
	`define ATCBMC300_M15S2 1'b1
`else
	`define ATCBMC300_M15S2 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV3
	`define ATCBMC300_M15S3 1'b1
`else
	`define ATCBMC300_M15S3 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV4
	`define ATCBMC300_M15S4 1'b1
`else
	`define ATCBMC300_M15S4 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV5
	`define ATCBMC300_M15S5 1'b1
`else
	`define ATCBMC300_M15S5 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV6
	`define ATCBMC300_M15S6 1'b1
`else
	`define ATCBMC300_M15S6 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV7
	`define ATCBMC300_M15S7 1'b1
`else
	`define ATCBMC300_M15S7 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV8
	`define ATCBMC300_M15S8 1'b1
`else
	`define ATCBMC300_M15S8 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV9
	`define ATCBMC300_M15S9 1'b1
`else
	`define ATCBMC300_M15S9 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV10
	`define ATCBMC300_M15S10 1'b1
`else
	`define ATCBMC300_M15S10 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV11
	`define ATCBMC300_M15S11 1'b1
`else
	`define ATCBMC300_M15S11 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV12
	`define ATCBMC300_M15S12 1'b1
`else
	`define ATCBMC300_M15S12 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV13
	`define ATCBMC300_M15S13 1'b1
`else
	`define ATCBMC300_M15S13 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV14
	`define ATCBMC300_M15S14 1'b1
`else
	`define ATCBMC300_M15S14 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV15
	`define ATCBMC300_M15S15 1'b1
`else
	`define ATCBMC300_M15S15 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV16
	`define ATCBMC300_M15S16 1'b1
`else
	`define ATCBMC300_M15S16 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV17
	`define ATCBMC300_M15S17 1'b1
`else
	`define ATCBMC300_M15S17 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV18
	`define ATCBMC300_M15S18 1'b1
`else
	`define ATCBMC300_M15S18 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV19
	`define ATCBMC300_M15S19 1'b1
`else
	`define ATCBMC300_M15S19 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV20
	`define ATCBMC300_M15S20 1'b1
`else
	`define ATCBMC300_M15S20 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV21
	`define ATCBMC300_M15S21 1'b1
`else
	`define ATCBMC300_M15S21 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV22
	`define ATCBMC300_M15S22 1'b1
`else
	`define ATCBMC300_M15S22 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV23
	`define ATCBMC300_M15S23 1'b1
`else
	`define ATCBMC300_M15S23 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV24
	`define ATCBMC300_M15S24 1'b1
`else
	`define ATCBMC300_M15S24 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV25
	`define ATCBMC300_M15S25 1'b1
`else
	`define ATCBMC300_M15S25 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV26
	`define ATCBMC300_M15S26 1'b1
`else
	`define ATCBMC300_M15S26 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV27
	`define ATCBMC300_M15S27 1'b1
`else
	`define ATCBMC300_M15S27 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV28
	`define ATCBMC300_M15S28 1'b1
`else
	`define ATCBMC300_M15S28 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV29
	`define ATCBMC300_M15S29 1'b1
`else
	`define ATCBMC300_M15S29 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV30
	`define ATCBMC300_M15S30 1'b1
`else
	`define ATCBMC300_M15S30 1'b0
`endif
`ifdef ATCBMC300_MST15_SLV31
	`define ATCBMC300_M15S31 1'b1
`else
	`define ATCBMC300_M15S31 1'b0
`endif
// VPERL_GENERATED_END
`endif
