
// This RTL design follows AE350P design spec V0.5.
//

module ae350_testgen (
// VPERL: &PORTLIST;
// VPERL_GENERATED_BEGIN
	  scan_test,
	  scan_enable 
// VPERL_GENERATED_END
);

output	scan_test;
output	scan_enable;


assign	scan_test	= 1'b0;
assign	scan_enable	= 1'b0;

endmodule
