`ifdef MACRO_CONVERTER_VH
`else
`define MACRO_CONVERTER_VH

// ATCBMC300_MxSx must have been defined in atcbmc300_const.vh. However,
// when random configuration is used, the content of atcbmc300_config.vh is
// not used so that all ATCBMC300_MxSx's are 1'b0. Override them when
// NDS_Mx_CONNS is defined. (At least one is defined).
//
// VPERL_BEGIN
// foreach $x (0 .. 15) {
//   :`ifdef NDS_M${x}_CONNS
//   foreach $y (0 .. 31) {
//     :	`undef ATCBMC300_M${x}S${y}
//     :	`define ATCBMC300_M${x}S${y}	(((`NDS_M${x}_CONNS>>$y) & 1) ? 1'b1 : 1'b0)
//   }
//   :`else	// !NDS_M${x}_CONNS
//   print "\t`define	NDS_M${x}_CONNS {";
//   for ($y = 31; $y > 0; $y--) {
//     print "`ATCBMC300_M${x}S${y}, ";
//   }
//   print "`ATCBMC300_M${x}S0}\n";
//   :`endif	// NDS_M${x}_CONNS
// }
// VPERL_END

// VPERL_GENERATED_BEGIN
`ifdef NDS_M0_CONNS
	`undef ATCBMC300_M0S0
	`define ATCBMC300_M0S0	(((`NDS_M0_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S1
	`define ATCBMC300_M0S1	(((`NDS_M0_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S2
	`define ATCBMC300_M0S2	(((`NDS_M0_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S3
	`define ATCBMC300_M0S3	(((`NDS_M0_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S4
	`define ATCBMC300_M0S4	(((`NDS_M0_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S5
	`define ATCBMC300_M0S5	(((`NDS_M0_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S6
	`define ATCBMC300_M0S6	(((`NDS_M0_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S7
	`define ATCBMC300_M0S7	(((`NDS_M0_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S8
	`define ATCBMC300_M0S8	(((`NDS_M0_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S9
	`define ATCBMC300_M0S9	(((`NDS_M0_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S10
	`define ATCBMC300_M0S10	(((`NDS_M0_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S11
	`define ATCBMC300_M0S11	(((`NDS_M0_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S12
	`define ATCBMC300_M0S12	(((`NDS_M0_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S13
	`define ATCBMC300_M0S13	(((`NDS_M0_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S14
	`define ATCBMC300_M0S14	(((`NDS_M0_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S15
	`define ATCBMC300_M0S15	(((`NDS_M0_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S16
	`define ATCBMC300_M0S16	(((`NDS_M0_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S17
	`define ATCBMC300_M0S17	(((`NDS_M0_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S18
	`define ATCBMC300_M0S18	(((`NDS_M0_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S19
	`define ATCBMC300_M0S19	(((`NDS_M0_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S20
	`define ATCBMC300_M0S20	(((`NDS_M0_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S21
	`define ATCBMC300_M0S21	(((`NDS_M0_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S22
	`define ATCBMC300_M0S22	(((`NDS_M0_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S23
	`define ATCBMC300_M0S23	(((`NDS_M0_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S24
	`define ATCBMC300_M0S24	(((`NDS_M0_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S25
	`define ATCBMC300_M0S25	(((`NDS_M0_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S26
	`define ATCBMC300_M0S26	(((`NDS_M0_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S27
	`define ATCBMC300_M0S27	(((`NDS_M0_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S28
	`define ATCBMC300_M0S28	(((`NDS_M0_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S29
	`define ATCBMC300_M0S29	(((`NDS_M0_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S30
	`define ATCBMC300_M0S30	(((`NDS_M0_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M0S31
	`define ATCBMC300_M0S31	(((`NDS_M0_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M0_CONNS
	`define	NDS_M0_CONNS {`ATCBMC300_M0S31, `ATCBMC300_M0S30, `ATCBMC300_M0S29, `ATCBMC300_M0S28, `ATCBMC300_M0S27, `ATCBMC300_M0S26, `ATCBMC300_M0S25, `ATCBMC300_M0S24, `ATCBMC300_M0S23, `ATCBMC300_M0S22, `ATCBMC300_M0S21, `ATCBMC300_M0S20, `ATCBMC300_M0S19, `ATCBMC300_M0S18, `ATCBMC300_M0S17, `ATCBMC300_M0S16, `ATCBMC300_M0S15, `ATCBMC300_M0S14, `ATCBMC300_M0S13, `ATCBMC300_M0S12, `ATCBMC300_M0S11, `ATCBMC300_M0S10, `ATCBMC300_M0S9, `ATCBMC300_M0S8, `ATCBMC300_M0S7, `ATCBMC300_M0S6, `ATCBMC300_M0S5, `ATCBMC300_M0S4, `ATCBMC300_M0S3, `ATCBMC300_M0S2, `ATCBMC300_M0S1, `ATCBMC300_M0S0}
`endif	// NDS_M0_CONNS
`ifdef NDS_M1_CONNS
	`undef ATCBMC300_M1S0
	`define ATCBMC300_M1S0	(((`NDS_M1_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S1
	`define ATCBMC300_M1S1	(((`NDS_M1_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S2
	`define ATCBMC300_M1S2	(((`NDS_M1_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S3
	`define ATCBMC300_M1S3	(((`NDS_M1_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S4
	`define ATCBMC300_M1S4	(((`NDS_M1_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S5
	`define ATCBMC300_M1S5	(((`NDS_M1_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S6
	`define ATCBMC300_M1S6	(((`NDS_M1_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S7
	`define ATCBMC300_M1S7	(((`NDS_M1_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S8
	`define ATCBMC300_M1S8	(((`NDS_M1_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S9
	`define ATCBMC300_M1S9	(((`NDS_M1_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S10
	`define ATCBMC300_M1S10	(((`NDS_M1_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S11
	`define ATCBMC300_M1S11	(((`NDS_M1_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S12
	`define ATCBMC300_M1S12	(((`NDS_M1_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S13
	`define ATCBMC300_M1S13	(((`NDS_M1_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S14
	`define ATCBMC300_M1S14	(((`NDS_M1_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S15
	`define ATCBMC300_M1S15	(((`NDS_M1_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S16
	`define ATCBMC300_M1S16	(((`NDS_M1_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S17
	`define ATCBMC300_M1S17	(((`NDS_M1_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S18
	`define ATCBMC300_M1S18	(((`NDS_M1_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S19
	`define ATCBMC300_M1S19	(((`NDS_M1_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S20
	`define ATCBMC300_M1S20	(((`NDS_M1_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S21
	`define ATCBMC300_M1S21	(((`NDS_M1_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S22
	`define ATCBMC300_M1S22	(((`NDS_M1_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S23
	`define ATCBMC300_M1S23	(((`NDS_M1_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S24
	`define ATCBMC300_M1S24	(((`NDS_M1_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S25
	`define ATCBMC300_M1S25	(((`NDS_M1_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S26
	`define ATCBMC300_M1S26	(((`NDS_M1_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S27
	`define ATCBMC300_M1S27	(((`NDS_M1_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S28
	`define ATCBMC300_M1S28	(((`NDS_M1_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S29
	`define ATCBMC300_M1S29	(((`NDS_M1_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S30
	`define ATCBMC300_M1S30	(((`NDS_M1_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M1S31
	`define ATCBMC300_M1S31	(((`NDS_M1_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M1_CONNS
	`define	NDS_M1_CONNS {`ATCBMC300_M1S31, `ATCBMC300_M1S30, `ATCBMC300_M1S29, `ATCBMC300_M1S28, `ATCBMC300_M1S27, `ATCBMC300_M1S26, `ATCBMC300_M1S25, `ATCBMC300_M1S24, `ATCBMC300_M1S23, `ATCBMC300_M1S22, `ATCBMC300_M1S21, `ATCBMC300_M1S20, `ATCBMC300_M1S19, `ATCBMC300_M1S18, `ATCBMC300_M1S17, `ATCBMC300_M1S16, `ATCBMC300_M1S15, `ATCBMC300_M1S14, `ATCBMC300_M1S13, `ATCBMC300_M1S12, `ATCBMC300_M1S11, `ATCBMC300_M1S10, `ATCBMC300_M1S9, `ATCBMC300_M1S8, `ATCBMC300_M1S7, `ATCBMC300_M1S6, `ATCBMC300_M1S5, `ATCBMC300_M1S4, `ATCBMC300_M1S3, `ATCBMC300_M1S2, `ATCBMC300_M1S1, `ATCBMC300_M1S0}
`endif	// NDS_M1_CONNS
`ifdef NDS_M2_CONNS
	`undef ATCBMC300_M2S0
	`define ATCBMC300_M2S0	(((`NDS_M2_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S1
	`define ATCBMC300_M2S1	(((`NDS_M2_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S2
	`define ATCBMC300_M2S2	(((`NDS_M2_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S3
	`define ATCBMC300_M2S3	(((`NDS_M2_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S4
	`define ATCBMC300_M2S4	(((`NDS_M2_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S5
	`define ATCBMC300_M2S5	(((`NDS_M2_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S6
	`define ATCBMC300_M2S6	(((`NDS_M2_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S7
	`define ATCBMC300_M2S7	(((`NDS_M2_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S8
	`define ATCBMC300_M2S8	(((`NDS_M2_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S9
	`define ATCBMC300_M2S9	(((`NDS_M2_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S10
	`define ATCBMC300_M2S10	(((`NDS_M2_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S11
	`define ATCBMC300_M2S11	(((`NDS_M2_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S12
	`define ATCBMC300_M2S12	(((`NDS_M2_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S13
	`define ATCBMC300_M2S13	(((`NDS_M2_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S14
	`define ATCBMC300_M2S14	(((`NDS_M2_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S15
	`define ATCBMC300_M2S15	(((`NDS_M2_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S16
	`define ATCBMC300_M2S16	(((`NDS_M2_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S17
	`define ATCBMC300_M2S17	(((`NDS_M2_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S18
	`define ATCBMC300_M2S18	(((`NDS_M2_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S19
	`define ATCBMC300_M2S19	(((`NDS_M2_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S20
	`define ATCBMC300_M2S20	(((`NDS_M2_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S21
	`define ATCBMC300_M2S21	(((`NDS_M2_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S22
	`define ATCBMC300_M2S22	(((`NDS_M2_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S23
	`define ATCBMC300_M2S23	(((`NDS_M2_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S24
	`define ATCBMC300_M2S24	(((`NDS_M2_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S25
	`define ATCBMC300_M2S25	(((`NDS_M2_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S26
	`define ATCBMC300_M2S26	(((`NDS_M2_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S27
	`define ATCBMC300_M2S27	(((`NDS_M2_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S28
	`define ATCBMC300_M2S28	(((`NDS_M2_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S29
	`define ATCBMC300_M2S29	(((`NDS_M2_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S30
	`define ATCBMC300_M2S30	(((`NDS_M2_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M2S31
	`define ATCBMC300_M2S31	(((`NDS_M2_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M2_CONNS
	`define	NDS_M2_CONNS {`ATCBMC300_M2S31, `ATCBMC300_M2S30, `ATCBMC300_M2S29, `ATCBMC300_M2S28, `ATCBMC300_M2S27, `ATCBMC300_M2S26, `ATCBMC300_M2S25, `ATCBMC300_M2S24, `ATCBMC300_M2S23, `ATCBMC300_M2S22, `ATCBMC300_M2S21, `ATCBMC300_M2S20, `ATCBMC300_M2S19, `ATCBMC300_M2S18, `ATCBMC300_M2S17, `ATCBMC300_M2S16, `ATCBMC300_M2S15, `ATCBMC300_M2S14, `ATCBMC300_M2S13, `ATCBMC300_M2S12, `ATCBMC300_M2S11, `ATCBMC300_M2S10, `ATCBMC300_M2S9, `ATCBMC300_M2S8, `ATCBMC300_M2S7, `ATCBMC300_M2S6, `ATCBMC300_M2S5, `ATCBMC300_M2S4, `ATCBMC300_M2S3, `ATCBMC300_M2S2, `ATCBMC300_M2S1, `ATCBMC300_M2S0}
`endif	// NDS_M2_CONNS
`ifdef NDS_M3_CONNS
	`undef ATCBMC300_M3S0
	`define ATCBMC300_M3S0	(((`NDS_M3_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S1
	`define ATCBMC300_M3S1	(((`NDS_M3_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S2
	`define ATCBMC300_M3S2	(((`NDS_M3_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S3
	`define ATCBMC300_M3S3	(((`NDS_M3_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S4
	`define ATCBMC300_M3S4	(((`NDS_M3_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S5
	`define ATCBMC300_M3S5	(((`NDS_M3_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S6
	`define ATCBMC300_M3S6	(((`NDS_M3_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S7
	`define ATCBMC300_M3S7	(((`NDS_M3_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S8
	`define ATCBMC300_M3S8	(((`NDS_M3_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S9
	`define ATCBMC300_M3S9	(((`NDS_M3_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S10
	`define ATCBMC300_M3S10	(((`NDS_M3_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S11
	`define ATCBMC300_M3S11	(((`NDS_M3_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S12
	`define ATCBMC300_M3S12	(((`NDS_M3_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S13
	`define ATCBMC300_M3S13	(((`NDS_M3_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S14
	`define ATCBMC300_M3S14	(((`NDS_M3_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S15
	`define ATCBMC300_M3S15	(((`NDS_M3_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S16
	`define ATCBMC300_M3S16	(((`NDS_M3_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S17
	`define ATCBMC300_M3S17	(((`NDS_M3_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S18
	`define ATCBMC300_M3S18	(((`NDS_M3_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S19
	`define ATCBMC300_M3S19	(((`NDS_M3_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S20
	`define ATCBMC300_M3S20	(((`NDS_M3_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S21
	`define ATCBMC300_M3S21	(((`NDS_M3_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S22
	`define ATCBMC300_M3S22	(((`NDS_M3_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S23
	`define ATCBMC300_M3S23	(((`NDS_M3_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S24
	`define ATCBMC300_M3S24	(((`NDS_M3_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S25
	`define ATCBMC300_M3S25	(((`NDS_M3_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S26
	`define ATCBMC300_M3S26	(((`NDS_M3_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S27
	`define ATCBMC300_M3S27	(((`NDS_M3_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S28
	`define ATCBMC300_M3S28	(((`NDS_M3_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S29
	`define ATCBMC300_M3S29	(((`NDS_M3_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S30
	`define ATCBMC300_M3S30	(((`NDS_M3_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M3S31
	`define ATCBMC300_M3S31	(((`NDS_M3_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M3_CONNS
	`define	NDS_M3_CONNS {`ATCBMC300_M3S31, `ATCBMC300_M3S30, `ATCBMC300_M3S29, `ATCBMC300_M3S28, `ATCBMC300_M3S27, `ATCBMC300_M3S26, `ATCBMC300_M3S25, `ATCBMC300_M3S24, `ATCBMC300_M3S23, `ATCBMC300_M3S22, `ATCBMC300_M3S21, `ATCBMC300_M3S20, `ATCBMC300_M3S19, `ATCBMC300_M3S18, `ATCBMC300_M3S17, `ATCBMC300_M3S16, `ATCBMC300_M3S15, `ATCBMC300_M3S14, `ATCBMC300_M3S13, `ATCBMC300_M3S12, `ATCBMC300_M3S11, `ATCBMC300_M3S10, `ATCBMC300_M3S9, `ATCBMC300_M3S8, `ATCBMC300_M3S7, `ATCBMC300_M3S6, `ATCBMC300_M3S5, `ATCBMC300_M3S4, `ATCBMC300_M3S3, `ATCBMC300_M3S2, `ATCBMC300_M3S1, `ATCBMC300_M3S0}
`endif	// NDS_M3_CONNS
`ifdef NDS_M4_CONNS
	`undef ATCBMC300_M4S0
	`define ATCBMC300_M4S0	(((`NDS_M4_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S1
	`define ATCBMC300_M4S1	(((`NDS_M4_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S2
	`define ATCBMC300_M4S2	(((`NDS_M4_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S3
	`define ATCBMC300_M4S3	(((`NDS_M4_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S4
	`define ATCBMC300_M4S4	(((`NDS_M4_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S5
	`define ATCBMC300_M4S5	(((`NDS_M4_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S6
	`define ATCBMC300_M4S6	(((`NDS_M4_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S7
	`define ATCBMC300_M4S7	(((`NDS_M4_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S8
	`define ATCBMC300_M4S8	(((`NDS_M4_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S9
	`define ATCBMC300_M4S9	(((`NDS_M4_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S10
	`define ATCBMC300_M4S10	(((`NDS_M4_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S11
	`define ATCBMC300_M4S11	(((`NDS_M4_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S12
	`define ATCBMC300_M4S12	(((`NDS_M4_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S13
	`define ATCBMC300_M4S13	(((`NDS_M4_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S14
	`define ATCBMC300_M4S14	(((`NDS_M4_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S15
	`define ATCBMC300_M4S15	(((`NDS_M4_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S16
	`define ATCBMC300_M4S16	(((`NDS_M4_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S17
	`define ATCBMC300_M4S17	(((`NDS_M4_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S18
	`define ATCBMC300_M4S18	(((`NDS_M4_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S19
	`define ATCBMC300_M4S19	(((`NDS_M4_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S20
	`define ATCBMC300_M4S20	(((`NDS_M4_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S21
	`define ATCBMC300_M4S21	(((`NDS_M4_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S22
	`define ATCBMC300_M4S22	(((`NDS_M4_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S23
	`define ATCBMC300_M4S23	(((`NDS_M4_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S24
	`define ATCBMC300_M4S24	(((`NDS_M4_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S25
	`define ATCBMC300_M4S25	(((`NDS_M4_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S26
	`define ATCBMC300_M4S26	(((`NDS_M4_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S27
	`define ATCBMC300_M4S27	(((`NDS_M4_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S28
	`define ATCBMC300_M4S28	(((`NDS_M4_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S29
	`define ATCBMC300_M4S29	(((`NDS_M4_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S30
	`define ATCBMC300_M4S30	(((`NDS_M4_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M4S31
	`define ATCBMC300_M4S31	(((`NDS_M4_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M4_CONNS
	`define	NDS_M4_CONNS {`ATCBMC300_M4S31, `ATCBMC300_M4S30, `ATCBMC300_M4S29, `ATCBMC300_M4S28, `ATCBMC300_M4S27, `ATCBMC300_M4S26, `ATCBMC300_M4S25, `ATCBMC300_M4S24, `ATCBMC300_M4S23, `ATCBMC300_M4S22, `ATCBMC300_M4S21, `ATCBMC300_M4S20, `ATCBMC300_M4S19, `ATCBMC300_M4S18, `ATCBMC300_M4S17, `ATCBMC300_M4S16, `ATCBMC300_M4S15, `ATCBMC300_M4S14, `ATCBMC300_M4S13, `ATCBMC300_M4S12, `ATCBMC300_M4S11, `ATCBMC300_M4S10, `ATCBMC300_M4S9, `ATCBMC300_M4S8, `ATCBMC300_M4S7, `ATCBMC300_M4S6, `ATCBMC300_M4S5, `ATCBMC300_M4S4, `ATCBMC300_M4S3, `ATCBMC300_M4S2, `ATCBMC300_M4S1, `ATCBMC300_M4S0}
`endif	// NDS_M4_CONNS
`ifdef NDS_M5_CONNS
	`undef ATCBMC300_M5S0
	`define ATCBMC300_M5S0	(((`NDS_M5_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S1
	`define ATCBMC300_M5S1	(((`NDS_M5_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S2
	`define ATCBMC300_M5S2	(((`NDS_M5_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S3
	`define ATCBMC300_M5S3	(((`NDS_M5_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S4
	`define ATCBMC300_M5S4	(((`NDS_M5_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S5
	`define ATCBMC300_M5S5	(((`NDS_M5_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S6
	`define ATCBMC300_M5S6	(((`NDS_M5_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S7
	`define ATCBMC300_M5S7	(((`NDS_M5_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S8
	`define ATCBMC300_M5S8	(((`NDS_M5_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S9
	`define ATCBMC300_M5S9	(((`NDS_M5_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S10
	`define ATCBMC300_M5S10	(((`NDS_M5_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S11
	`define ATCBMC300_M5S11	(((`NDS_M5_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S12
	`define ATCBMC300_M5S12	(((`NDS_M5_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S13
	`define ATCBMC300_M5S13	(((`NDS_M5_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S14
	`define ATCBMC300_M5S14	(((`NDS_M5_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S15
	`define ATCBMC300_M5S15	(((`NDS_M5_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S16
	`define ATCBMC300_M5S16	(((`NDS_M5_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S17
	`define ATCBMC300_M5S17	(((`NDS_M5_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S18
	`define ATCBMC300_M5S18	(((`NDS_M5_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S19
	`define ATCBMC300_M5S19	(((`NDS_M5_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S20
	`define ATCBMC300_M5S20	(((`NDS_M5_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S21
	`define ATCBMC300_M5S21	(((`NDS_M5_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S22
	`define ATCBMC300_M5S22	(((`NDS_M5_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S23
	`define ATCBMC300_M5S23	(((`NDS_M5_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S24
	`define ATCBMC300_M5S24	(((`NDS_M5_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S25
	`define ATCBMC300_M5S25	(((`NDS_M5_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S26
	`define ATCBMC300_M5S26	(((`NDS_M5_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S27
	`define ATCBMC300_M5S27	(((`NDS_M5_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S28
	`define ATCBMC300_M5S28	(((`NDS_M5_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S29
	`define ATCBMC300_M5S29	(((`NDS_M5_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S30
	`define ATCBMC300_M5S30	(((`NDS_M5_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M5S31
	`define ATCBMC300_M5S31	(((`NDS_M5_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M5_CONNS
	`define	NDS_M5_CONNS {`ATCBMC300_M5S31, `ATCBMC300_M5S30, `ATCBMC300_M5S29, `ATCBMC300_M5S28, `ATCBMC300_M5S27, `ATCBMC300_M5S26, `ATCBMC300_M5S25, `ATCBMC300_M5S24, `ATCBMC300_M5S23, `ATCBMC300_M5S22, `ATCBMC300_M5S21, `ATCBMC300_M5S20, `ATCBMC300_M5S19, `ATCBMC300_M5S18, `ATCBMC300_M5S17, `ATCBMC300_M5S16, `ATCBMC300_M5S15, `ATCBMC300_M5S14, `ATCBMC300_M5S13, `ATCBMC300_M5S12, `ATCBMC300_M5S11, `ATCBMC300_M5S10, `ATCBMC300_M5S9, `ATCBMC300_M5S8, `ATCBMC300_M5S7, `ATCBMC300_M5S6, `ATCBMC300_M5S5, `ATCBMC300_M5S4, `ATCBMC300_M5S3, `ATCBMC300_M5S2, `ATCBMC300_M5S1, `ATCBMC300_M5S0}
`endif	// NDS_M5_CONNS
`ifdef NDS_M6_CONNS
	`undef ATCBMC300_M6S0
	`define ATCBMC300_M6S0	(((`NDS_M6_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S1
	`define ATCBMC300_M6S1	(((`NDS_M6_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S2
	`define ATCBMC300_M6S2	(((`NDS_M6_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S3
	`define ATCBMC300_M6S3	(((`NDS_M6_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S4
	`define ATCBMC300_M6S4	(((`NDS_M6_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S5
	`define ATCBMC300_M6S5	(((`NDS_M6_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S6
	`define ATCBMC300_M6S6	(((`NDS_M6_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S7
	`define ATCBMC300_M6S7	(((`NDS_M6_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S8
	`define ATCBMC300_M6S8	(((`NDS_M6_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S9
	`define ATCBMC300_M6S9	(((`NDS_M6_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S10
	`define ATCBMC300_M6S10	(((`NDS_M6_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S11
	`define ATCBMC300_M6S11	(((`NDS_M6_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S12
	`define ATCBMC300_M6S12	(((`NDS_M6_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S13
	`define ATCBMC300_M6S13	(((`NDS_M6_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S14
	`define ATCBMC300_M6S14	(((`NDS_M6_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S15
	`define ATCBMC300_M6S15	(((`NDS_M6_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S16
	`define ATCBMC300_M6S16	(((`NDS_M6_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S17
	`define ATCBMC300_M6S17	(((`NDS_M6_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S18
	`define ATCBMC300_M6S18	(((`NDS_M6_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S19
	`define ATCBMC300_M6S19	(((`NDS_M6_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S20
	`define ATCBMC300_M6S20	(((`NDS_M6_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S21
	`define ATCBMC300_M6S21	(((`NDS_M6_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S22
	`define ATCBMC300_M6S22	(((`NDS_M6_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S23
	`define ATCBMC300_M6S23	(((`NDS_M6_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S24
	`define ATCBMC300_M6S24	(((`NDS_M6_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S25
	`define ATCBMC300_M6S25	(((`NDS_M6_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S26
	`define ATCBMC300_M6S26	(((`NDS_M6_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S27
	`define ATCBMC300_M6S27	(((`NDS_M6_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S28
	`define ATCBMC300_M6S28	(((`NDS_M6_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S29
	`define ATCBMC300_M6S29	(((`NDS_M6_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S30
	`define ATCBMC300_M6S30	(((`NDS_M6_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M6S31
	`define ATCBMC300_M6S31	(((`NDS_M6_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M6_CONNS
	`define	NDS_M6_CONNS {`ATCBMC300_M6S31, `ATCBMC300_M6S30, `ATCBMC300_M6S29, `ATCBMC300_M6S28, `ATCBMC300_M6S27, `ATCBMC300_M6S26, `ATCBMC300_M6S25, `ATCBMC300_M6S24, `ATCBMC300_M6S23, `ATCBMC300_M6S22, `ATCBMC300_M6S21, `ATCBMC300_M6S20, `ATCBMC300_M6S19, `ATCBMC300_M6S18, `ATCBMC300_M6S17, `ATCBMC300_M6S16, `ATCBMC300_M6S15, `ATCBMC300_M6S14, `ATCBMC300_M6S13, `ATCBMC300_M6S12, `ATCBMC300_M6S11, `ATCBMC300_M6S10, `ATCBMC300_M6S9, `ATCBMC300_M6S8, `ATCBMC300_M6S7, `ATCBMC300_M6S6, `ATCBMC300_M6S5, `ATCBMC300_M6S4, `ATCBMC300_M6S3, `ATCBMC300_M6S2, `ATCBMC300_M6S1, `ATCBMC300_M6S0}
`endif	// NDS_M6_CONNS
`ifdef NDS_M7_CONNS
	`undef ATCBMC300_M7S0
	`define ATCBMC300_M7S0	(((`NDS_M7_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S1
	`define ATCBMC300_M7S1	(((`NDS_M7_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S2
	`define ATCBMC300_M7S2	(((`NDS_M7_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S3
	`define ATCBMC300_M7S3	(((`NDS_M7_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S4
	`define ATCBMC300_M7S4	(((`NDS_M7_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S5
	`define ATCBMC300_M7S5	(((`NDS_M7_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S6
	`define ATCBMC300_M7S6	(((`NDS_M7_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S7
	`define ATCBMC300_M7S7	(((`NDS_M7_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S8
	`define ATCBMC300_M7S8	(((`NDS_M7_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S9
	`define ATCBMC300_M7S9	(((`NDS_M7_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S10
	`define ATCBMC300_M7S10	(((`NDS_M7_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S11
	`define ATCBMC300_M7S11	(((`NDS_M7_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S12
	`define ATCBMC300_M7S12	(((`NDS_M7_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S13
	`define ATCBMC300_M7S13	(((`NDS_M7_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S14
	`define ATCBMC300_M7S14	(((`NDS_M7_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S15
	`define ATCBMC300_M7S15	(((`NDS_M7_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S16
	`define ATCBMC300_M7S16	(((`NDS_M7_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S17
	`define ATCBMC300_M7S17	(((`NDS_M7_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S18
	`define ATCBMC300_M7S18	(((`NDS_M7_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S19
	`define ATCBMC300_M7S19	(((`NDS_M7_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S20
	`define ATCBMC300_M7S20	(((`NDS_M7_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S21
	`define ATCBMC300_M7S21	(((`NDS_M7_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S22
	`define ATCBMC300_M7S22	(((`NDS_M7_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S23
	`define ATCBMC300_M7S23	(((`NDS_M7_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S24
	`define ATCBMC300_M7S24	(((`NDS_M7_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S25
	`define ATCBMC300_M7S25	(((`NDS_M7_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S26
	`define ATCBMC300_M7S26	(((`NDS_M7_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S27
	`define ATCBMC300_M7S27	(((`NDS_M7_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S28
	`define ATCBMC300_M7S28	(((`NDS_M7_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S29
	`define ATCBMC300_M7S29	(((`NDS_M7_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S30
	`define ATCBMC300_M7S30	(((`NDS_M7_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M7S31
	`define ATCBMC300_M7S31	(((`NDS_M7_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M7_CONNS
	`define	NDS_M7_CONNS {`ATCBMC300_M7S31, `ATCBMC300_M7S30, `ATCBMC300_M7S29, `ATCBMC300_M7S28, `ATCBMC300_M7S27, `ATCBMC300_M7S26, `ATCBMC300_M7S25, `ATCBMC300_M7S24, `ATCBMC300_M7S23, `ATCBMC300_M7S22, `ATCBMC300_M7S21, `ATCBMC300_M7S20, `ATCBMC300_M7S19, `ATCBMC300_M7S18, `ATCBMC300_M7S17, `ATCBMC300_M7S16, `ATCBMC300_M7S15, `ATCBMC300_M7S14, `ATCBMC300_M7S13, `ATCBMC300_M7S12, `ATCBMC300_M7S11, `ATCBMC300_M7S10, `ATCBMC300_M7S9, `ATCBMC300_M7S8, `ATCBMC300_M7S7, `ATCBMC300_M7S6, `ATCBMC300_M7S5, `ATCBMC300_M7S4, `ATCBMC300_M7S3, `ATCBMC300_M7S2, `ATCBMC300_M7S1, `ATCBMC300_M7S0}
`endif	// NDS_M7_CONNS
`ifdef NDS_M8_CONNS
	`undef ATCBMC300_M8S0
	`define ATCBMC300_M8S0	(((`NDS_M8_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S1
	`define ATCBMC300_M8S1	(((`NDS_M8_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S2
	`define ATCBMC300_M8S2	(((`NDS_M8_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S3
	`define ATCBMC300_M8S3	(((`NDS_M8_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S4
	`define ATCBMC300_M8S4	(((`NDS_M8_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S5
	`define ATCBMC300_M8S5	(((`NDS_M8_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S6
	`define ATCBMC300_M8S6	(((`NDS_M8_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S7
	`define ATCBMC300_M8S7	(((`NDS_M8_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S8
	`define ATCBMC300_M8S8	(((`NDS_M8_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S9
	`define ATCBMC300_M8S9	(((`NDS_M8_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S10
	`define ATCBMC300_M8S10	(((`NDS_M8_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S11
	`define ATCBMC300_M8S11	(((`NDS_M8_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S12
	`define ATCBMC300_M8S12	(((`NDS_M8_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S13
	`define ATCBMC300_M8S13	(((`NDS_M8_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S14
	`define ATCBMC300_M8S14	(((`NDS_M8_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S15
	`define ATCBMC300_M8S15	(((`NDS_M8_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S16
	`define ATCBMC300_M8S16	(((`NDS_M8_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S17
	`define ATCBMC300_M8S17	(((`NDS_M8_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S18
	`define ATCBMC300_M8S18	(((`NDS_M8_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S19
	`define ATCBMC300_M8S19	(((`NDS_M8_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S20
	`define ATCBMC300_M8S20	(((`NDS_M8_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S21
	`define ATCBMC300_M8S21	(((`NDS_M8_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S22
	`define ATCBMC300_M8S22	(((`NDS_M8_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S23
	`define ATCBMC300_M8S23	(((`NDS_M8_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S24
	`define ATCBMC300_M8S24	(((`NDS_M8_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S25
	`define ATCBMC300_M8S25	(((`NDS_M8_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S26
	`define ATCBMC300_M8S26	(((`NDS_M8_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S27
	`define ATCBMC300_M8S27	(((`NDS_M8_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S28
	`define ATCBMC300_M8S28	(((`NDS_M8_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S29
	`define ATCBMC300_M8S29	(((`NDS_M8_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S30
	`define ATCBMC300_M8S30	(((`NDS_M8_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M8S31
	`define ATCBMC300_M8S31	(((`NDS_M8_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M8_CONNS
	`define	NDS_M8_CONNS {`ATCBMC300_M8S31, `ATCBMC300_M8S30, `ATCBMC300_M8S29, `ATCBMC300_M8S28, `ATCBMC300_M8S27, `ATCBMC300_M8S26, `ATCBMC300_M8S25, `ATCBMC300_M8S24, `ATCBMC300_M8S23, `ATCBMC300_M8S22, `ATCBMC300_M8S21, `ATCBMC300_M8S20, `ATCBMC300_M8S19, `ATCBMC300_M8S18, `ATCBMC300_M8S17, `ATCBMC300_M8S16, `ATCBMC300_M8S15, `ATCBMC300_M8S14, `ATCBMC300_M8S13, `ATCBMC300_M8S12, `ATCBMC300_M8S11, `ATCBMC300_M8S10, `ATCBMC300_M8S9, `ATCBMC300_M8S8, `ATCBMC300_M8S7, `ATCBMC300_M8S6, `ATCBMC300_M8S5, `ATCBMC300_M8S4, `ATCBMC300_M8S3, `ATCBMC300_M8S2, `ATCBMC300_M8S1, `ATCBMC300_M8S0}
`endif	// NDS_M8_CONNS
`ifdef NDS_M9_CONNS
	`undef ATCBMC300_M9S0
	`define ATCBMC300_M9S0	(((`NDS_M9_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S1
	`define ATCBMC300_M9S1	(((`NDS_M9_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S2
	`define ATCBMC300_M9S2	(((`NDS_M9_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S3
	`define ATCBMC300_M9S3	(((`NDS_M9_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S4
	`define ATCBMC300_M9S4	(((`NDS_M9_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S5
	`define ATCBMC300_M9S5	(((`NDS_M9_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S6
	`define ATCBMC300_M9S6	(((`NDS_M9_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S7
	`define ATCBMC300_M9S7	(((`NDS_M9_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S8
	`define ATCBMC300_M9S8	(((`NDS_M9_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S9
	`define ATCBMC300_M9S9	(((`NDS_M9_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S10
	`define ATCBMC300_M9S10	(((`NDS_M9_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S11
	`define ATCBMC300_M9S11	(((`NDS_M9_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S12
	`define ATCBMC300_M9S12	(((`NDS_M9_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S13
	`define ATCBMC300_M9S13	(((`NDS_M9_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S14
	`define ATCBMC300_M9S14	(((`NDS_M9_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S15
	`define ATCBMC300_M9S15	(((`NDS_M9_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S16
	`define ATCBMC300_M9S16	(((`NDS_M9_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S17
	`define ATCBMC300_M9S17	(((`NDS_M9_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S18
	`define ATCBMC300_M9S18	(((`NDS_M9_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S19
	`define ATCBMC300_M9S19	(((`NDS_M9_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S20
	`define ATCBMC300_M9S20	(((`NDS_M9_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S21
	`define ATCBMC300_M9S21	(((`NDS_M9_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S22
	`define ATCBMC300_M9S22	(((`NDS_M9_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S23
	`define ATCBMC300_M9S23	(((`NDS_M9_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S24
	`define ATCBMC300_M9S24	(((`NDS_M9_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S25
	`define ATCBMC300_M9S25	(((`NDS_M9_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S26
	`define ATCBMC300_M9S26	(((`NDS_M9_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S27
	`define ATCBMC300_M9S27	(((`NDS_M9_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S28
	`define ATCBMC300_M9S28	(((`NDS_M9_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S29
	`define ATCBMC300_M9S29	(((`NDS_M9_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S30
	`define ATCBMC300_M9S30	(((`NDS_M9_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M9S31
	`define ATCBMC300_M9S31	(((`NDS_M9_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M9_CONNS
	`define	NDS_M9_CONNS {`ATCBMC300_M9S31, `ATCBMC300_M9S30, `ATCBMC300_M9S29, `ATCBMC300_M9S28, `ATCBMC300_M9S27, `ATCBMC300_M9S26, `ATCBMC300_M9S25, `ATCBMC300_M9S24, `ATCBMC300_M9S23, `ATCBMC300_M9S22, `ATCBMC300_M9S21, `ATCBMC300_M9S20, `ATCBMC300_M9S19, `ATCBMC300_M9S18, `ATCBMC300_M9S17, `ATCBMC300_M9S16, `ATCBMC300_M9S15, `ATCBMC300_M9S14, `ATCBMC300_M9S13, `ATCBMC300_M9S12, `ATCBMC300_M9S11, `ATCBMC300_M9S10, `ATCBMC300_M9S9, `ATCBMC300_M9S8, `ATCBMC300_M9S7, `ATCBMC300_M9S6, `ATCBMC300_M9S5, `ATCBMC300_M9S4, `ATCBMC300_M9S3, `ATCBMC300_M9S2, `ATCBMC300_M9S1, `ATCBMC300_M9S0}
`endif	// NDS_M9_CONNS
`ifdef NDS_M10_CONNS
	`undef ATCBMC300_M10S0
	`define ATCBMC300_M10S0	(((`NDS_M10_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S1
	`define ATCBMC300_M10S1	(((`NDS_M10_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S2
	`define ATCBMC300_M10S2	(((`NDS_M10_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S3
	`define ATCBMC300_M10S3	(((`NDS_M10_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S4
	`define ATCBMC300_M10S4	(((`NDS_M10_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S5
	`define ATCBMC300_M10S5	(((`NDS_M10_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S6
	`define ATCBMC300_M10S6	(((`NDS_M10_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S7
	`define ATCBMC300_M10S7	(((`NDS_M10_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S8
	`define ATCBMC300_M10S8	(((`NDS_M10_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S9
	`define ATCBMC300_M10S9	(((`NDS_M10_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S10
	`define ATCBMC300_M10S10	(((`NDS_M10_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S11
	`define ATCBMC300_M10S11	(((`NDS_M10_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S12
	`define ATCBMC300_M10S12	(((`NDS_M10_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S13
	`define ATCBMC300_M10S13	(((`NDS_M10_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S14
	`define ATCBMC300_M10S14	(((`NDS_M10_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S15
	`define ATCBMC300_M10S15	(((`NDS_M10_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S16
	`define ATCBMC300_M10S16	(((`NDS_M10_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S17
	`define ATCBMC300_M10S17	(((`NDS_M10_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S18
	`define ATCBMC300_M10S18	(((`NDS_M10_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S19
	`define ATCBMC300_M10S19	(((`NDS_M10_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S20
	`define ATCBMC300_M10S20	(((`NDS_M10_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S21
	`define ATCBMC300_M10S21	(((`NDS_M10_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S22
	`define ATCBMC300_M10S22	(((`NDS_M10_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S23
	`define ATCBMC300_M10S23	(((`NDS_M10_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S24
	`define ATCBMC300_M10S24	(((`NDS_M10_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S25
	`define ATCBMC300_M10S25	(((`NDS_M10_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S26
	`define ATCBMC300_M10S26	(((`NDS_M10_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S27
	`define ATCBMC300_M10S27	(((`NDS_M10_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S28
	`define ATCBMC300_M10S28	(((`NDS_M10_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S29
	`define ATCBMC300_M10S29	(((`NDS_M10_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S30
	`define ATCBMC300_M10S30	(((`NDS_M10_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M10S31
	`define ATCBMC300_M10S31	(((`NDS_M10_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M10_CONNS
	`define	NDS_M10_CONNS {`ATCBMC300_M10S31, `ATCBMC300_M10S30, `ATCBMC300_M10S29, `ATCBMC300_M10S28, `ATCBMC300_M10S27, `ATCBMC300_M10S26, `ATCBMC300_M10S25, `ATCBMC300_M10S24, `ATCBMC300_M10S23, `ATCBMC300_M10S22, `ATCBMC300_M10S21, `ATCBMC300_M10S20, `ATCBMC300_M10S19, `ATCBMC300_M10S18, `ATCBMC300_M10S17, `ATCBMC300_M10S16, `ATCBMC300_M10S15, `ATCBMC300_M10S14, `ATCBMC300_M10S13, `ATCBMC300_M10S12, `ATCBMC300_M10S11, `ATCBMC300_M10S10, `ATCBMC300_M10S9, `ATCBMC300_M10S8, `ATCBMC300_M10S7, `ATCBMC300_M10S6, `ATCBMC300_M10S5, `ATCBMC300_M10S4, `ATCBMC300_M10S3, `ATCBMC300_M10S2, `ATCBMC300_M10S1, `ATCBMC300_M10S0}
`endif	// NDS_M10_CONNS
`ifdef NDS_M11_CONNS
	`undef ATCBMC300_M11S0
	`define ATCBMC300_M11S0	(((`NDS_M11_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S1
	`define ATCBMC300_M11S1	(((`NDS_M11_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S2
	`define ATCBMC300_M11S2	(((`NDS_M11_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S3
	`define ATCBMC300_M11S3	(((`NDS_M11_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S4
	`define ATCBMC300_M11S4	(((`NDS_M11_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S5
	`define ATCBMC300_M11S5	(((`NDS_M11_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S6
	`define ATCBMC300_M11S6	(((`NDS_M11_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S7
	`define ATCBMC300_M11S7	(((`NDS_M11_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S8
	`define ATCBMC300_M11S8	(((`NDS_M11_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S9
	`define ATCBMC300_M11S9	(((`NDS_M11_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S10
	`define ATCBMC300_M11S10	(((`NDS_M11_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S11
	`define ATCBMC300_M11S11	(((`NDS_M11_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S12
	`define ATCBMC300_M11S12	(((`NDS_M11_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S13
	`define ATCBMC300_M11S13	(((`NDS_M11_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S14
	`define ATCBMC300_M11S14	(((`NDS_M11_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S15
	`define ATCBMC300_M11S15	(((`NDS_M11_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S16
	`define ATCBMC300_M11S16	(((`NDS_M11_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S17
	`define ATCBMC300_M11S17	(((`NDS_M11_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S18
	`define ATCBMC300_M11S18	(((`NDS_M11_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S19
	`define ATCBMC300_M11S19	(((`NDS_M11_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S20
	`define ATCBMC300_M11S20	(((`NDS_M11_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S21
	`define ATCBMC300_M11S21	(((`NDS_M11_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S22
	`define ATCBMC300_M11S22	(((`NDS_M11_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S23
	`define ATCBMC300_M11S23	(((`NDS_M11_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S24
	`define ATCBMC300_M11S24	(((`NDS_M11_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S25
	`define ATCBMC300_M11S25	(((`NDS_M11_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S26
	`define ATCBMC300_M11S26	(((`NDS_M11_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S27
	`define ATCBMC300_M11S27	(((`NDS_M11_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S28
	`define ATCBMC300_M11S28	(((`NDS_M11_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S29
	`define ATCBMC300_M11S29	(((`NDS_M11_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S30
	`define ATCBMC300_M11S30	(((`NDS_M11_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M11S31
	`define ATCBMC300_M11S31	(((`NDS_M11_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M11_CONNS
	`define	NDS_M11_CONNS {`ATCBMC300_M11S31, `ATCBMC300_M11S30, `ATCBMC300_M11S29, `ATCBMC300_M11S28, `ATCBMC300_M11S27, `ATCBMC300_M11S26, `ATCBMC300_M11S25, `ATCBMC300_M11S24, `ATCBMC300_M11S23, `ATCBMC300_M11S22, `ATCBMC300_M11S21, `ATCBMC300_M11S20, `ATCBMC300_M11S19, `ATCBMC300_M11S18, `ATCBMC300_M11S17, `ATCBMC300_M11S16, `ATCBMC300_M11S15, `ATCBMC300_M11S14, `ATCBMC300_M11S13, `ATCBMC300_M11S12, `ATCBMC300_M11S11, `ATCBMC300_M11S10, `ATCBMC300_M11S9, `ATCBMC300_M11S8, `ATCBMC300_M11S7, `ATCBMC300_M11S6, `ATCBMC300_M11S5, `ATCBMC300_M11S4, `ATCBMC300_M11S3, `ATCBMC300_M11S2, `ATCBMC300_M11S1, `ATCBMC300_M11S0}
`endif	// NDS_M11_CONNS
`ifdef NDS_M12_CONNS
	`undef ATCBMC300_M12S0
	`define ATCBMC300_M12S0	(((`NDS_M12_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S1
	`define ATCBMC300_M12S1	(((`NDS_M12_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S2
	`define ATCBMC300_M12S2	(((`NDS_M12_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S3
	`define ATCBMC300_M12S3	(((`NDS_M12_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S4
	`define ATCBMC300_M12S4	(((`NDS_M12_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S5
	`define ATCBMC300_M12S5	(((`NDS_M12_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S6
	`define ATCBMC300_M12S6	(((`NDS_M12_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S7
	`define ATCBMC300_M12S7	(((`NDS_M12_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S8
	`define ATCBMC300_M12S8	(((`NDS_M12_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S9
	`define ATCBMC300_M12S9	(((`NDS_M12_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S10
	`define ATCBMC300_M12S10	(((`NDS_M12_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S11
	`define ATCBMC300_M12S11	(((`NDS_M12_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S12
	`define ATCBMC300_M12S12	(((`NDS_M12_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S13
	`define ATCBMC300_M12S13	(((`NDS_M12_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S14
	`define ATCBMC300_M12S14	(((`NDS_M12_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S15
	`define ATCBMC300_M12S15	(((`NDS_M12_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S16
	`define ATCBMC300_M12S16	(((`NDS_M12_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S17
	`define ATCBMC300_M12S17	(((`NDS_M12_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S18
	`define ATCBMC300_M12S18	(((`NDS_M12_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S19
	`define ATCBMC300_M12S19	(((`NDS_M12_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S20
	`define ATCBMC300_M12S20	(((`NDS_M12_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S21
	`define ATCBMC300_M12S21	(((`NDS_M12_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S22
	`define ATCBMC300_M12S22	(((`NDS_M12_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S23
	`define ATCBMC300_M12S23	(((`NDS_M12_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S24
	`define ATCBMC300_M12S24	(((`NDS_M12_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S25
	`define ATCBMC300_M12S25	(((`NDS_M12_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S26
	`define ATCBMC300_M12S26	(((`NDS_M12_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S27
	`define ATCBMC300_M12S27	(((`NDS_M12_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S28
	`define ATCBMC300_M12S28	(((`NDS_M12_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S29
	`define ATCBMC300_M12S29	(((`NDS_M12_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S30
	`define ATCBMC300_M12S30	(((`NDS_M12_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M12S31
	`define ATCBMC300_M12S31	(((`NDS_M12_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M12_CONNS
	`define	NDS_M12_CONNS {`ATCBMC300_M12S31, `ATCBMC300_M12S30, `ATCBMC300_M12S29, `ATCBMC300_M12S28, `ATCBMC300_M12S27, `ATCBMC300_M12S26, `ATCBMC300_M12S25, `ATCBMC300_M12S24, `ATCBMC300_M12S23, `ATCBMC300_M12S22, `ATCBMC300_M12S21, `ATCBMC300_M12S20, `ATCBMC300_M12S19, `ATCBMC300_M12S18, `ATCBMC300_M12S17, `ATCBMC300_M12S16, `ATCBMC300_M12S15, `ATCBMC300_M12S14, `ATCBMC300_M12S13, `ATCBMC300_M12S12, `ATCBMC300_M12S11, `ATCBMC300_M12S10, `ATCBMC300_M12S9, `ATCBMC300_M12S8, `ATCBMC300_M12S7, `ATCBMC300_M12S6, `ATCBMC300_M12S5, `ATCBMC300_M12S4, `ATCBMC300_M12S3, `ATCBMC300_M12S2, `ATCBMC300_M12S1, `ATCBMC300_M12S0}
`endif	// NDS_M12_CONNS
`ifdef NDS_M13_CONNS
	`undef ATCBMC300_M13S0
	`define ATCBMC300_M13S0	(((`NDS_M13_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S1
	`define ATCBMC300_M13S1	(((`NDS_M13_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S2
	`define ATCBMC300_M13S2	(((`NDS_M13_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S3
	`define ATCBMC300_M13S3	(((`NDS_M13_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S4
	`define ATCBMC300_M13S4	(((`NDS_M13_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S5
	`define ATCBMC300_M13S5	(((`NDS_M13_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S6
	`define ATCBMC300_M13S6	(((`NDS_M13_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S7
	`define ATCBMC300_M13S7	(((`NDS_M13_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S8
	`define ATCBMC300_M13S8	(((`NDS_M13_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S9
	`define ATCBMC300_M13S9	(((`NDS_M13_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S10
	`define ATCBMC300_M13S10	(((`NDS_M13_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S11
	`define ATCBMC300_M13S11	(((`NDS_M13_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S12
	`define ATCBMC300_M13S12	(((`NDS_M13_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S13
	`define ATCBMC300_M13S13	(((`NDS_M13_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S14
	`define ATCBMC300_M13S14	(((`NDS_M13_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S15
	`define ATCBMC300_M13S15	(((`NDS_M13_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S16
	`define ATCBMC300_M13S16	(((`NDS_M13_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S17
	`define ATCBMC300_M13S17	(((`NDS_M13_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S18
	`define ATCBMC300_M13S18	(((`NDS_M13_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S19
	`define ATCBMC300_M13S19	(((`NDS_M13_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S20
	`define ATCBMC300_M13S20	(((`NDS_M13_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S21
	`define ATCBMC300_M13S21	(((`NDS_M13_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S22
	`define ATCBMC300_M13S22	(((`NDS_M13_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S23
	`define ATCBMC300_M13S23	(((`NDS_M13_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S24
	`define ATCBMC300_M13S24	(((`NDS_M13_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S25
	`define ATCBMC300_M13S25	(((`NDS_M13_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S26
	`define ATCBMC300_M13S26	(((`NDS_M13_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S27
	`define ATCBMC300_M13S27	(((`NDS_M13_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S28
	`define ATCBMC300_M13S28	(((`NDS_M13_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S29
	`define ATCBMC300_M13S29	(((`NDS_M13_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S30
	`define ATCBMC300_M13S30	(((`NDS_M13_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M13S31
	`define ATCBMC300_M13S31	(((`NDS_M13_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M13_CONNS
	`define	NDS_M13_CONNS {`ATCBMC300_M13S31, `ATCBMC300_M13S30, `ATCBMC300_M13S29, `ATCBMC300_M13S28, `ATCBMC300_M13S27, `ATCBMC300_M13S26, `ATCBMC300_M13S25, `ATCBMC300_M13S24, `ATCBMC300_M13S23, `ATCBMC300_M13S22, `ATCBMC300_M13S21, `ATCBMC300_M13S20, `ATCBMC300_M13S19, `ATCBMC300_M13S18, `ATCBMC300_M13S17, `ATCBMC300_M13S16, `ATCBMC300_M13S15, `ATCBMC300_M13S14, `ATCBMC300_M13S13, `ATCBMC300_M13S12, `ATCBMC300_M13S11, `ATCBMC300_M13S10, `ATCBMC300_M13S9, `ATCBMC300_M13S8, `ATCBMC300_M13S7, `ATCBMC300_M13S6, `ATCBMC300_M13S5, `ATCBMC300_M13S4, `ATCBMC300_M13S3, `ATCBMC300_M13S2, `ATCBMC300_M13S1, `ATCBMC300_M13S0}
`endif	// NDS_M13_CONNS
`ifdef NDS_M14_CONNS
	`undef ATCBMC300_M14S0
	`define ATCBMC300_M14S0	(((`NDS_M14_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S1
	`define ATCBMC300_M14S1	(((`NDS_M14_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S2
	`define ATCBMC300_M14S2	(((`NDS_M14_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S3
	`define ATCBMC300_M14S3	(((`NDS_M14_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S4
	`define ATCBMC300_M14S4	(((`NDS_M14_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S5
	`define ATCBMC300_M14S5	(((`NDS_M14_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S6
	`define ATCBMC300_M14S6	(((`NDS_M14_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S7
	`define ATCBMC300_M14S7	(((`NDS_M14_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S8
	`define ATCBMC300_M14S8	(((`NDS_M14_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S9
	`define ATCBMC300_M14S9	(((`NDS_M14_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S10
	`define ATCBMC300_M14S10	(((`NDS_M14_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S11
	`define ATCBMC300_M14S11	(((`NDS_M14_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S12
	`define ATCBMC300_M14S12	(((`NDS_M14_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S13
	`define ATCBMC300_M14S13	(((`NDS_M14_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S14
	`define ATCBMC300_M14S14	(((`NDS_M14_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S15
	`define ATCBMC300_M14S15	(((`NDS_M14_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S16
	`define ATCBMC300_M14S16	(((`NDS_M14_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S17
	`define ATCBMC300_M14S17	(((`NDS_M14_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S18
	`define ATCBMC300_M14S18	(((`NDS_M14_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S19
	`define ATCBMC300_M14S19	(((`NDS_M14_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S20
	`define ATCBMC300_M14S20	(((`NDS_M14_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S21
	`define ATCBMC300_M14S21	(((`NDS_M14_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S22
	`define ATCBMC300_M14S22	(((`NDS_M14_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S23
	`define ATCBMC300_M14S23	(((`NDS_M14_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S24
	`define ATCBMC300_M14S24	(((`NDS_M14_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S25
	`define ATCBMC300_M14S25	(((`NDS_M14_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S26
	`define ATCBMC300_M14S26	(((`NDS_M14_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S27
	`define ATCBMC300_M14S27	(((`NDS_M14_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S28
	`define ATCBMC300_M14S28	(((`NDS_M14_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S29
	`define ATCBMC300_M14S29	(((`NDS_M14_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S30
	`define ATCBMC300_M14S30	(((`NDS_M14_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M14S31
	`define ATCBMC300_M14S31	(((`NDS_M14_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M14_CONNS
	`define	NDS_M14_CONNS {`ATCBMC300_M14S31, `ATCBMC300_M14S30, `ATCBMC300_M14S29, `ATCBMC300_M14S28, `ATCBMC300_M14S27, `ATCBMC300_M14S26, `ATCBMC300_M14S25, `ATCBMC300_M14S24, `ATCBMC300_M14S23, `ATCBMC300_M14S22, `ATCBMC300_M14S21, `ATCBMC300_M14S20, `ATCBMC300_M14S19, `ATCBMC300_M14S18, `ATCBMC300_M14S17, `ATCBMC300_M14S16, `ATCBMC300_M14S15, `ATCBMC300_M14S14, `ATCBMC300_M14S13, `ATCBMC300_M14S12, `ATCBMC300_M14S11, `ATCBMC300_M14S10, `ATCBMC300_M14S9, `ATCBMC300_M14S8, `ATCBMC300_M14S7, `ATCBMC300_M14S6, `ATCBMC300_M14S5, `ATCBMC300_M14S4, `ATCBMC300_M14S3, `ATCBMC300_M14S2, `ATCBMC300_M14S1, `ATCBMC300_M14S0}
`endif	// NDS_M14_CONNS
`ifdef NDS_M15_CONNS
	`undef ATCBMC300_M15S0
	`define ATCBMC300_M15S0	(((`NDS_M15_CONNS>>0) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S1
	`define ATCBMC300_M15S1	(((`NDS_M15_CONNS>>1) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S2
	`define ATCBMC300_M15S2	(((`NDS_M15_CONNS>>2) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S3
	`define ATCBMC300_M15S3	(((`NDS_M15_CONNS>>3) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S4
	`define ATCBMC300_M15S4	(((`NDS_M15_CONNS>>4) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S5
	`define ATCBMC300_M15S5	(((`NDS_M15_CONNS>>5) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S6
	`define ATCBMC300_M15S6	(((`NDS_M15_CONNS>>6) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S7
	`define ATCBMC300_M15S7	(((`NDS_M15_CONNS>>7) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S8
	`define ATCBMC300_M15S8	(((`NDS_M15_CONNS>>8) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S9
	`define ATCBMC300_M15S9	(((`NDS_M15_CONNS>>9) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S10
	`define ATCBMC300_M15S10	(((`NDS_M15_CONNS>>10) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S11
	`define ATCBMC300_M15S11	(((`NDS_M15_CONNS>>11) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S12
	`define ATCBMC300_M15S12	(((`NDS_M15_CONNS>>12) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S13
	`define ATCBMC300_M15S13	(((`NDS_M15_CONNS>>13) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S14
	`define ATCBMC300_M15S14	(((`NDS_M15_CONNS>>14) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S15
	`define ATCBMC300_M15S15	(((`NDS_M15_CONNS>>15) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S16
	`define ATCBMC300_M15S16	(((`NDS_M15_CONNS>>16) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S17
	`define ATCBMC300_M15S17	(((`NDS_M15_CONNS>>17) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S18
	`define ATCBMC300_M15S18	(((`NDS_M15_CONNS>>18) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S19
	`define ATCBMC300_M15S19	(((`NDS_M15_CONNS>>19) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S20
	`define ATCBMC300_M15S20	(((`NDS_M15_CONNS>>20) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S21
	`define ATCBMC300_M15S21	(((`NDS_M15_CONNS>>21) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S22
	`define ATCBMC300_M15S22	(((`NDS_M15_CONNS>>22) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S23
	`define ATCBMC300_M15S23	(((`NDS_M15_CONNS>>23) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S24
	`define ATCBMC300_M15S24	(((`NDS_M15_CONNS>>24) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S25
	`define ATCBMC300_M15S25	(((`NDS_M15_CONNS>>25) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S26
	`define ATCBMC300_M15S26	(((`NDS_M15_CONNS>>26) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S27
	`define ATCBMC300_M15S27	(((`NDS_M15_CONNS>>27) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S28
	`define ATCBMC300_M15S28	(((`NDS_M15_CONNS>>28) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S29
	`define ATCBMC300_M15S29	(((`NDS_M15_CONNS>>29) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S30
	`define ATCBMC300_M15S30	(((`NDS_M15_CONNS>>30) & 1) ? 1'b1 : 1'b0)
	`undef ATCBMC300_M15S31
	`define ATCBMC300_M15S31	(((`NDS_M15_CONNS>>31) & 1) ? 1'b1 : 1'b0)
`else	// !NDS_M15_CONNS
	`define	NDS_M15_CONNS {`ATCBMC300_M15S31, `ATCBMC300_M15S30, `ATCBMC300_M15S29, `ATCBMC300_M15S28, `ATCBMC300_M15S27, `ATCBMC300_M15S26, `ATCBMC300_M15S25, `ATCBMC300_M15S24, `ATCBMC300_M15S23, `ATCBMC300_M15S22, `ATCBMC300_M15S21, `ATCBMC300_M15S20, `ATCBMC300_M15S19, `ATCBMC300_M15S18, `ATCBMC300_M15S17, `ATCBMC300_M15S16, `ATCBMC300_M15S15, `ATCBMC300_M15S14, `ATCBMC300_M15S13, `ATCBMC300_M15S12, `ATCBMC300_M15S11, `ATCBMC300_M15S10, `ATCBMC300_M15S9, `ATCBMC300_M15S8, `ATCBMC300_M15S7, `ATCBMC300_M15S6, `ATCBMC300_M15S5, `ATCBMC300_M15S4, `ATCBMC300_M15S3, `ATCBMC300_M15S2, `ATCBMC300_M15S1, `ATCBMC300_M15S0}
`endif	// NDS_M15_CONNS
// VPERL_GENERATED_END
`endif
