`timescale 1ns/1ps
`include "xmr.vh"

`include "atcbmc300_config.vh"
`include "atcbmc300_const.vh"

`ifdef NDS_AXI_MASTER_MODEL_PAT
	`ifdef WITH_COV		// Block coverage.
		`define NDS_COV_ENABLED		// Used in axi_master.pat.
	`elsif WITH_EXP_COV	// Expression coverage.
		`define NDS_COV_ENABLED		// Used in axi_master.pat.
	`endif
`endif	// NDS_AXI_MASTER_MODEL_PAT

`ifndef ATCBMC300_ADDR_WIDTH
	`define ATCBMC300_ADDR_WIDTH		32
`endif

`ifndef ATCBMC300_ID_WIDTH
	`define ATCBMC300_ID_WIDTH		4
`endif

`ifndef NDS_ERROR_PROBABILITY
	`define NDS_ERROR_PROBABILITY		10		// %.
`endif

`ifndef NDS_DEFAULT_DELAY_MAX
	`define NDS_DEFAULT_DELAY_MAX		10		// Cycles.
`endif

`ifndef NDS_DEFAULT_TRANS_NUM
	`define NDS_DEFAULT_TRANS_NUM		500		// Transaction#.
`endif

// For the performance, disable errors.
`ifdef NDS_PERFORMANCE_TEST
	`undef NDS_ERROR_PROBABILITY
	`define NDS_ERROR_PROBABILITY		0

	`undef NDS_DEFAULT_DELAY_MAX
	`define NDS_DEFAULT_DELAY_MAX		0

	// VPERL_BEGIN
	// for $x (0 .. 15) {
	//   :`ifdef NDS_MST${x}_DELAY_MAX
	//   :	`undef NDS_MST${x}_DELAY_MAX
	//   :`endif
	// }
	// VPERL_END

	// VPERL_GENERATED_BEGIN
	`ifdef NDS_MST0_DELAY_MAX
		`undef NDS_MST0_DELAY_MAX
	`endif
	`ifdef NDS_MST1_DELAY_MAX
		`undef NDS_MST1_DELAY_MAX
	`endif
	`ifdef NDS_MST2_DELAY_MAX
		`undef NDS_MST2_DELAY_MAX
	`endif
	`ifdef NDS_MST3_DELAY_MAX
		`undef NDS_MST3_DELAY_MAX
	`endif
	`ifdef NDS_MST4_DELAY_MAX
		`undef NDS_MST4_DELAY_MAX
	`endif
	`ifdef NDS_MST5_DELAY_MAX
		`undef NDS_MST5_DELAY_MAX
	`endif
	`ifdef NDS_MST6_DELAY_MAX
		`undef NDS_MST6_DELAY_MAX
	`endif
	`ifdef NDS_MST7_DELAY_MAX
		`undef NDS_MST7_DELAY_MAX
	`endif
	`ifdef NDS_MST8_DELAY_MAX
		`undef NDS_MST8_DELAY_MAX
	`endif
	`ifdef NDS_MST9_DELAY_MAX
		`undef NDS_MST9_DELAY_MAX
	`endif
	`ifdef NDS_MST10_DELAY_MAX
		`undef NDS_MST10_DELAY_MAX
	`endif
	`ifdef NDS_MST11_DELAY_MAX
		`undef NDS_MST11_DELAY_MAX
	`endif
	`ifdef NDS_MST12_DELAY_MAX
		`undef NDS_MST12_DELAY_MAX
	`endif
	`ifdef NDS_MST13_DELAY_MAX
		`undef NDS_MST13_DELAY_MAX
	`endif
	`ifdef NDS_MST14_DELAY_MAX
		`undef NDS_MST14_DELAY_MAX
	`endif
	`ifdef NDS_MST15_DELAY_MAX
		`undef NDS_MST15_DELAY_MAX
	`endif
	// VPERL_GENERATED_END
`endif

// Translate macros.
`include "macro_convert.vh"

package cfg_pkg;	// Config package.
	parameter unsigned	MID_WIDTH = 8;		// Model ID width (Not AXI's).
	parameter unsigned	US_ID_WIDTH = `ATCBMC300_ID_WIDTH;	// Master's AXI ID width.
	parameter unsigned	DS_ID_WIDTH = `ATCBMC300_ID_WIDTH+4;	// Slave's AXI ID width.

	typedef logic [MID_WIDTH-1:0]	mid_t;
	typedef logic [US_ID_WIDTH-1:0]	us_id_t;
	typedef logic [DS_ID_WIDTH-1:0]	ds_id_t;
endpackage: cfg_pkg

// VPERL_BEGIN
// 
// &MODULE("system");
//
// ### Configurable parameters ###
//
// &PARAM("ADDR_WIDTH = `ATCBMC300_ADDR_WIDTH");
//
// ### Derived or fixed parameters ###
//
// &PARAM("DATA_BYTES = `ATCBMC300_DATA_WIDTH / 8");
// &PARAM("DATA_SIZE = \$clog2(DATA_BYTES)");
// &PARAM("DATA_WIDTH = 8 * DATA_BYTES");
// &PARAM("DATA_MSB = DATA_WIDTH - 1");
// &PARAM("US_ID_WIDTH = `ATCBMC300_ID_WIDTH");
// &PARAM("DS_ID_WIDTH = `ATCBMC300_ID_WIDTH+4");
//
// # ==========
// # DUT
// # ==========
// &INSTANCE("$PVC_LOCALDIR/andes_ip/peripheral_ip/atcbmc300/hdl/atcbmc300.v", "bmc300", {
// });
// &CONNECT("bmc300", {
// });
//
// # ==========
// # tb & model
// # ==========
// &INSTANCE("$PVC_LOCALDIR/andes_ip/peripheral_ip/atcbmc300/bench/blk_tb.sv", "bench", {
//	ADDR_WIDTH		=> "ADDR_WIDTH",
//	DATA_SIZE		=> "DATA_SIZE",
//	ERROR_PROBABILITY	=> "`NDS_ERROR_PROBABILITY",
//	DS_ID_WIDTH		=> "DS_ID_WIDTH",
// });
//
// foreach $i (0 .. 15) {
//   &IFDEF("ATCBMC300_MST${i}_SUPPORT");
//
//   &FORCE("wire", "us${i}_arlock");
//   &FORCE("wire", "us${i}_awlock");
//   &INSTANCE("$PVC_LOCALDIR/andes_vip/models/axi/hdl/axi_master_model.sv", "axi_master${i}", {
//      ADDR_WIDTH	=> "ADDR_WIDTH",
//   	DATA_WIDTH	=> "DATA_SIZE",
//   	ADDR_START	=> "0",
//      ADDR_SIZE	=> "(1<<ADDR_WIDTH)",
//   	MODEL_ID	=> ${i},
//	ID_WIDTH	=> "US_ID_WIDTH",
//	AXI4		=> "1'b1",
//	AXI4_AXLEN_LT16	=> "1'b0",
//	UNALIGN_SUPPORT	=> "1'b1",
//	MAX_BUF_DEPTH	=> 256,
//	WAIT_TIMEOUT_CNT=> 1000000,
//	DELAY_MAX	=> "`ifdef NDS_MST${i}_DELAY_MAX `NDS_MST${i}_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif",
//	TRANS_NUM	=> "`ifdef NDS_MST${i}_TRANS_NUM `NDS_MST${i}_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif",
//   });
//   &CONNECT("axi_master${i}", {
//     arvalid		=> "us${i}_arvalid",
//     arready		=> "us${i}_arready",
//     arburst		=> "us${i}_arburst",
//     arsize		=> "us${i}_arsize",
//     arlen		=> "us${i}_arlen",
//     araddr		=> "us${i}_araddr",
//     arid		=> "us${i}_arid",
//     arcache		=> "us${i}_arcache",
//     arlock		=> "{us${i}_arlock_b1, us${i}_arlock}",
//     arprot		=> "us${i}_arprot",
//     awvalid		=> "us${i}_awvalid",
//     awready		=> "us${i}_awready",
//     awburst		=> "us${i}_awburst",
//     awsize		=> "us${i}_awsize",
//     awlen		=> "us${i}_awlen",
//     awaddr		=> "us${i}_awaddr",
//     awid		=> "us${i}_awid",
//     awcache		=> "us${i}_awcache",
//     awlock		=> "{us${i}_awlock_b1, us${i}_awlock}",
//     awprot		=> "us${i}_awprot",
//     bvalid		=> "us${i}_bvalid",
//     bready		=> "us${i}_bready",
//     bid		=> "us${i}_bid",
//     bresp		=> "us${i}_bresp",
//     rvalid		=> "us${i}_rvalid",
//     rready		=> "us${i}_rready",
//     rid		=> "us${i}_rid",
//     rresp		=> "us${i}_rresp",
//     rlast		=> "us${i}_rlast",
//     rdata		=> "us${i}_rdata",
//     wvalid		=> "us${i}_wvalid",
//     wready		=> "us${i}_wready",
//     wid		=> "us${i}_wid",
//     wlast		=> "us${i}_wlast",
//     wstrb		=> "us${i}_wstrb",
//     wdata		=> "us${i}_wdata",
//   });
//
//   &INSTANCE("$PVC_LOCALDIR/andes_vip/monitors/hdl/axi_monitor.v", "axi_monitor_m${i}", {
//      ADDR_WIDTH	=> "ADDR_WIDTH",
//   	DATA_WIDTH	=> "DATA_SIZE",
//   	ID_WIDTH	=> "US_ID_WIDTH",
//   	MASTER_ID	=> ${i},
//   	SLAVE_ID	=> ${i},
//   	AXI4		=> "1'b1",
//   });
//   &CONNECT("axi_monitor_m${i}", {
//     arvalid		=> "us${i}_arvalid",
//     arready		=> "us${i}_arready",
//     arburst		=> "us${i}_arburst",
//     arsize		=> "us${i}_arsize",
//     arlen		=> "us${i}_arlen",
//     araddr		=> "us${i}_araddr",
//     arid		=> "us${i}_arid",
//     arcache		=> "us${i}_arcache",
//     arlock		=> "{us${i}_arlock_b1, us${i}_arlock}",
//     arprot		=> "us${i}_arprot",
//     awvalid		=> "us${i}_awvalid",
//     awready		=> "us${i}_awready",
//     awburst		=> "us${i}_awburst",
//     awsize		=> "us${i}_awsize",
//     awlen		=> "us${i}_awlen",
//     awaddr		=> "us${i}_awaddr",
//     awid		=> "us${i}_awid",
//     awcache		=> "us${i}_awcache",
//     awlock		=> "{us${i}_awlock_b1, us${i}_awlock}",
//     awprot		=> "us${i}_awprot",
//     bvalid		=> "us${i}_bvalid",
//     bready		=> "us${i}_bready",
//     bid		=> "us${i}_bid",
//     bresp		=> "us${i}_bresp",
//     rvalid		=> "us${i}_rvalid",
//     rready		=> "us${i}_rready",
//     rid		=> "us${i}_rid",
//     rresp		=> "us${i}_rresp",
//     rlast		=> "us${i}_rlast",
//     rdata		=> "us${i}_rdata",
//     wvalid		=> "us${i}_wvalid",
//     wready		=> "us${i}_wready",
//     wid		=> "us${i}_wid",
//     wlast		=> "us${i}_wlast",
//     wstrb		=> "us${i}_wstrb",
//     wdata		=> "us${i}_wdata",
//   });
//
//   &ENDIF();
// }
//
// foreach $i (1 .. 31) {
//   &IFDEF("ATCBMC300_SLV${i}_SUPPORT");
//
//   &INSTANCE("$PVC_LOCALDIR/andes_vip/models/axi/hdl/axi_slave_model.v", "axi_slave${i}", {
//     ADDR_WIDTH	=> "ADDR_WIDTH",
//     DATA_WIDTH	=> "DATA_SIZE",
//     ID_WIDTH		=> "DS_ID_WIDTH",
//     MEM_ADDR_WIDTH	=> "`ATCBMC300_SLV${i}_SIZE+19",
//     ADDR_DECODE_WIDTH=> "`ATCBMC300_SLV${i}_SIZE+19",
//     AXI4		=> "1'b1",
//     RAND_INIT_ON_READ_X	=> "1'b1",
//   });
//   &CONNECT("axi_slave${i}", {
//     arvalid		=> "ds${i}_arvalid",
//     arready		=> "ds${i}_arready",
//     arburst		=> "ds${i}_arburst",
//     arsize		=> "ds${i}_arsize",
//     arlen		=> "ds${i}_arlen",
//     araddr		=> "ds${i}_araddr",
//     arid		=> "ds${i}_arid",
//     arcache		=> "ds${i}_arcache",
//     arlock		=> "{1'b0, ds${i}_arlock}",
//     arprot		=> "ds${i}_arprot",
//     awvalid		=> "ds${i}_awvalid",
//     awready		=> "ds${i}_awready",
//     awburst		=> "ds${i}_awburst",
//     awsize		=> "ds${i}_awsize",
//     awlen		=> "ds${i}_awlen",
//     awaddr		=> "ds${i}_awaddr",
//     awid		=> "ds${i}_awid",
//     awcache		=> "ds${i}_awcache",
//     awlock		=> "{1'b0, ds${i}_awlock}",
//     awprot		=> "ds${i}_awprot",
//     bvalid		=> "ds${i}_bvalid",
//     bready		=> "ds${i}_bready",
//     bid		=> "ds${i}_bid",
//     bresp		=> "ds${i}_bresp",
//     rvalid		=> "ds${i}_rvalid",
//     rready		=> "ds${i}_rready",
//     rid		=> "ds${i}_rid",
//     rresp		=> "ds${i}_rresp",
//     rlast		=> "ds${i}_rlast",
//     rdata		=> "ds${i}_rdata",
//     wvalid		=> "ds${i}_wvalid",
//     wready		=> "ds${i}_wready",
//     wid		=> "ds${i}_wid",
//     wlast		=> "ds${i}_wlast",
//     wstrb		=> "ds${i}_wstrb",
//     wdata		=> "ds${i}_wdata",
//     csysreq		=> "1'b0",
//     csysack		=> "",
//     cactive		=> "",
//   });
//   &FORCE("supply0", "ds${i}_wid[DS_ID_WIDTH-1:0]");
//
//   &INSTANCE("$PVC_LOCALDIR/andes_vip/monitors/hdl/axi_monitor.v", "axi_monitor_s${i}", {
//     ADDR_WIDTH	=> "ADDR_WIDTH",
//     DATA_WIDTH	=> "DATA_SIZE",
//     ID_WIDTH		=> "DS_ID_WIDTH",
//     MASTER_ID	=> 100+${i},
//     SLAVE_ID		=> 100+${i},
//     AXI4		=> "1'b1",
//   });
//   &CONNECT("axi_monitor_s${i}", {
//     arvalid		=> "ds${i}_arvalid",
//     arready		=> "ds${i}_arready",
//     arburst		=> "ds${i}_arburst",
//     arsize		=> "ds${i}_arsize",
//     arlen		=> "ds${i}_arlen",
//     araddr		=> "ds${i}_araddr",
//     arid		=> "ds${i}_arid",
//     arcache		=> "ds${i}_arcache",
//     arlock		=> "{1'b0, ds${i}_arlock}",
//     arprot		=> "ds${i}_arprot",
//     awvalid		=> "ds${i}_awvalid",
//     awready		=> "ds${i}_awready",
//     awburst		=> "ds${i}_awburst",
//     awsize		=> "ds${i}_awsize",
//     awlen		=> "ds${i}_awlen",
//     awaddr		=> "ds${i}_awaddr",
//     awid		=> "ds${i}_awid",
//     awcache		=> "ds${i}_awcache",
//     awlock		=> "{1'b0, ds${i}_awlock}",
//     awprot		=> "ds${i}_awprot",
//     bvalid		=> "ds${i}_bvalid",
//     bready		=> "ds${i}_bready",
//     bid		=> "ds${i}_bid",
//     bresp		=> "ds${i}_bresp",
//     rvalid		=> "ds${i}_rvalid",
//     rready		=> "ds${i}_rready",
//     rid		=> "ds${i}_rid",
//     rresp		=> "ds${i}_rresp",
//     rlast		=> "ds${i}_rlast",
//     rdata		=> "ds${i}_rdata",
//     wvalid		=> "ds${i}_wvalid",
//     wready		=> "ds${i}_wready",
//     wid		=> "ds${i}_wid",
//     wlast		=> "ds${i}_wlast",
//     wstrb		=> "ds${i}_wstrb",
//     wdata		=> "ds${i}_wdata",
//   });
//
//   &ENDIF();
// }
//
// : `ifdef NDS_SCOREBOARD_EN
// : // scoreboard
// : blk_scb  blk_scb();
// :
// foreach $i (0 .. 15) {
// : `ifdef ATCBMC300_MST${i}_SUPPORT
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.SCB_ID_WIDTH = 8;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.AXI4 = 1'b1;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.CAPTURE_LOCK = 1'b1;
// : defparam `NDS_SYSTEM.axi_master${i}.scb_axim_mon.CAPTURE_ID = 1'b1;
// : `endif
// }
// :
// foreach $i (1 .. 31) {
// : `ifdef ATCBMC300_SLV${i}_SUPPORT
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.SCB_ID_WIDTH = 8;
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.AXI4 = 1'b1;
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.CAPTURE_LOCK = 1'b1;
// : defparam `NDS_SYSTEM.axi_slave${i}.scb_axis_mon.CAPTURE_ID = 1'b1;
// : `ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
// : defparam `NDS_SYSTEM.axi_slave${i}.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
// : `endif
// : `endif
// }
// : `endif // NDS_SCOREBOARD_EN
// :
//
// &ENDMODULE;
// : `ifdef NDS_SCOREBOARD_EN
// foreach $i (0 .. 15) {
// : `ifdef ATCBMC300_MST${i}_SUPPORT
// : bind axi_master_model :`NDS_SYSTEM.axi_master${i} scb_axim_mon scb_axim_mon (.*, .model_id(8'd${i}));
// : `endif
// }
// :
// foreach $i (1 .. 31) {
// : `ifdef ATCBMC300_SLV${i}_SUPPORT
// : bind axi_slave_model : `NDS_SYSTEM.axi_slave${i} scb_axis_mon scb_axis_mon (.*, .model_id(8'd${i}));
// : `endif
// }
// : `endif // NDS_SCOREBOARD_EN
//
// VPERL_END

// VPERL_GENERATED_BEGIN
module system (
);

parameter ADDR_WIDTH = `ATCBMC300_ADDR_WIDTH;
parameter DATA_BYTES = `ATCBMC300_DATA_WIDTH / 8;
parameter DATA_SIZE = $clog2(DATA_BYTES);
parameter DATA_WIDTH = 8 * DATA_BYTES;
parameter DATA_MSB = DATA_WIDTH - 1;
parameter US_ID_WIDTH = `ATCBMC300_ID_WIDTH;
parameter DS_ID_WIDTH = `ATCBMC300_ID_WIDTH+4;
`ifdef ATCBMC300_MST0_SUPPORT
wire                               [ADDR_WIDTH-1:0] us0_araddr;
wire                                          [1:0] us0_arburst;
wire                                          [3:0] us0_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us0_arid;
wire                                          [7:0] us0_arlen;
wire                                                us0_arlock;
wire                                                us0_arlock_b1;
wire                                          [2:0] us0_arprot;
wire                                          [2:0] us0_arsize;
wire                                                us0_arvalid;
wire                               [ADDR_WIDTH-1:0] us0_awaddr;
wire                                          [1:0] us0_awburst;
wire                                          [3:0] us0_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us0_awid;
wire                                          [7:0] us0_awlen;
wire                                                us0_awlock;
wire                                                us0_awlock_b1;
wire                                          [2:0] us0_awprot;
wire                                          [2:0] us0_awsize;
wire                                                us0_awvalid;
wire                                                us0_bready;
wire                                                us0_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us0_wdata;
wire                              [US_ID_WIDTH-1:0] us0_wid;
wire                                                us0_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us0_wstrb;
wire                                                us0_wvalid;
wire                                                us0_arready;
wire                                                us0_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us0_bid;
wire                                          [1:0] us0_bresp;
wire                                                us0_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us0_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us0_rid;
wire                                                us0_rlast;
wire                                          [1:0] us0_rresp;
wire                                                us0_rvalid;
wire                                                us0_wready;
`endif // ATCBMC300_MST0_SUPPORT
`ifdef ATCBMC300_SLV1_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds1_wid;
wire                                                ds1_arready;
wire                                                ds1_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds1_bid;
wire                                          [1:0] ds1_bresp;
wire                                                ds1_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds1_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds1_rid;
wire                                                ds1_rlast;
wire                                          [1:0] ds1_rresp;
wire                                                ds1_rvalid;
wire                                                ds1_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds1_araddr;
wire                                          [1:0] ds1_arburst;
wire                                          [3:0] ds1_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds1_arid;
wire                                          [7:0] ds1_arlen;
wire                                                ds1_arlock;
wire                                          [2:0] ds1_arprot;
wire                                          [2:0] ds1_arsize;
wire                                                ds1_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds1_awaddr;
wire                                          [1:0] ds1_awburst;
wire                                          [3:0] ds1_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds1_awid;
wire                                          [7:0] ds1_awlen;
wire                                                ds1_awlock;
wire                                          [2:0] ds1_awprot;
wire                                          [2:0] ds1_awsize;
wire                                                ds1_awvalid;
wire                                                ds1_bready;
wire                                                ds1_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds1_wdata;
wire                                                ds1_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds1_wstrb;
wire                                                ds1_wvalid;
`endif // ATCBMC300_SLV1_SUPPORT
`ifdef ATCBMC300_SLV2_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds2_wid;
wire                                                ds2_arready;
wire                                                ds2_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds2_bid;
wire                                          [1:0] ds2_bresp;
wire                                                ds2_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds2_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds2_rid;
wire                                                ds2_rlast;
wire                                          [1:0] ds2_rresp;
wire                                                ds2_rvalid;
wire                                                ds2_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds2_araddr;
wire                                          [1:0] ds2_arburst;
wire                                          [3:0] ds2_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds2_arid;
wire                                          [7:0] ds2_arlen;
wire                                                ds2_arlock;
wire                                          [2:0] ds2_arprot;
wire                                          [2:0] ds2_arsize;
wire                                                ds2_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds2_awaddr;
wire                                          [1:0] ds2_awburst;
wire                                          [3:0] ds2_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds2_awid;
wire                                          [7:0] ds2_awlen;
wire                                                ds2_awlock;
wire                                          [2:0] ds2_awprot;
wire                                          [2:0] ds2_awsize;
wire                                                ds2_awvalid;
wire                                                ds2_bready;
wire                                                ds2_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds2_wdata;
wire                                                ds2_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds2_wstrb;
wire                                                ds2_wvalid;
`endif // ATCBMC300_SLV2_SUPPORT
`ifdef ATCBMC300_SLV3_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds3_wid;
wire                                                ds3_arready;
wire                                                ds3_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds3_bid;
wire                                          [1:0] ds3_bresp;
wire                                                ds3_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds3_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds3_rid;
wire                                                ds3_rlast;
wire                                          [1:0] ds3_rresp;
wire                                                ds3_rvalid;
wire                                                ds3_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds3_araddr;
wire                                          [1:0] ds3_arburst;
wire                                          [3:0] ds3_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds3_arid;
wire                                          [7:0] ds3_arlen;
wire                                                ds3_arlock;
wire                                          [2:0] ds3_arprot;
wire                                          [2:0] ds3_arsize;
wire                                                ds3_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds3_awaddr;
wire                                          [1:0] ds3_awburst;
wire                                          [3:0] ds3_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds3_awid;
wire                                          [7:0] ds3_awlen;
wire                                                ds3_awlock;
wire                                          [2:0] ds3_awprot;
wire                                          [2:0] ds3_awsize;
wire                                                ds3_awvalid;
wire                                                ds3_bready;
wire                                                ds3_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds3_wdata;
wire                                                ds3_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds3_wstrb;
wire                                                ds3_wvalid;
`endif // ATCBMC300_SLV3_SUPPORT
`ifdef ATCBMC300_SLV4_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds4_wid;
wire                                                ds4_arready;
wire                                                ds4_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds4_bid;
wire                                          [1:0] ds4_bresp;
wire                                                ds4_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds4_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds4_rid;
wire                                                ds4_rlast;
wire                                          [1:0] ds4_rresp;
wire                                                ds4_rvalid;
wire                                                ds4_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds4_araddr;
wire                                          [1:0] ds4_arburst;
wire                                          [3:0] ds4_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds4_arid;
wire                                          [7:0] ds4_arlen;
wire                                                ds4_arlock;
wire                                          [2:0] ds4_arprot;
wire                                          [2:0] ds4_arsize;
wire                                                ds4_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds4_awaddr;
wire                                          [1:0] ds4_awburst;
wire                                          [3:0] ds4_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds4_awid;
wire                                          [7:0] ds4_awlen;
wire                                                ds4_awlock;
wire                                          [2:0] ds4_awprot;
wire                                          [2:0] ds4_awsize;
wire                                                ds4_awvalid;
wire                                                ds4_bready;
wire                                                ds4_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds4_wdata;
wire                                                ds4_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds4_wstrb;
wire                                                ds4_wvalid;
`endif // ATCBMC300_SLV4_SUPPORT
`ifdef ATCBMC300_SLV5_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds5_wid;
wire                                                ds5_arready;
wire                                                ds5_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds5_bid;
wire                                          [1:0] ds5_bresp;
wire                                                ds5_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds5_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds5_rid;
wire                                                ds5_rlast;
wire                                          [1:0] ds5_rresp;
wire                                                ds5_rvalid;
wire                                                ds5_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds5_araddr;
wire                                          [1:0] ds5_arburst;
wire                                          [3:0] ds5_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds5_arid;
wire                                          [7:0] ds5_arlen;
wire                                                ds5_arlock;
wire                                          [2:0] ds5_arprot;
wire                                          [2:0] ds5_arsize;
wire                                                ds5_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds5_awaddr;
wire                                          [1:0] ds5_awburst;
wire                                          [3:0] ds5_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds5_awid;
wire                                          [7:0] ds5_awlen;
wire                                                ds5_awlock;
wire                                          [2:0] ds5_awprot;
wire                                          [2:0] ds5_awsize;
wire                                                ds5_awvalid;
wire                                                ds5_bready;
wire                                                ds5_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds5_wdata;
wire                                                ds5_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds5_wstrb;
wire                                                ds5_wvalid;
`endif // ATCBMC300_SLV5_SUPPORT
`ifdef ATCBMC300_SLV6_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds6_wid;
wire                                                ds6_arready;
wire                                                ds6_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds6_bid;
wire                                          [1:0] ds6_bresp;
wire                                                ds6_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds6_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds6_rid;
wire                                                ds6_rlast;
wire                                          [1:0] ds6_rresp;
wire                                                ds6_rvalid;
wire                                                ds6_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds6_araddr;
wire                                          [1:0] ds6_arburst;
wire                                          [3:0] ds6_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds6_arid;
wire                                          [7:0] ds6_arlen;
wire                                                ds6_arlock;
wire                                          [2:0] ds6_arprot;
wire                                          [2:0] ds6_arsize;
wire                                                ds6_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds6_awaddr;
wire                                          [1:0] ds6_awburst;
wire                                          [3:0] ds6_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds6_awid;
wire                                          [7:0] ds6_awlen;
wire                                                ds6_awlock;
wire                                          [2:0] ds6_awprot;
wire                                          [2:0] ds6_awsize;
wire                                                ds6_awvalid;
wire                                                ds6_bready;
wire                                                ds6_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds6_wdata;
wire                                                ds6_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds6_wstrb;
wire                                                ds6_wvalid;
`endif // ATCBMC300_SLV6_SUPPORT
`ifdef ATCBMC300_SLV7_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds7_wid;
wire                                                ds7_arready;
wire                                                ds7_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds7_bid;
wire                                          [1:0] ds7_bresp;
wire                                                ds7_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds7_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds7_rid;
wire                                                ds7_rlast;
wire                                          [1:0] ds7_rresp;
wire                                                ds7_rvalid;
wire                                                ds7_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds7_araddr;
wire                                          [1:0] ds7_arburst;
wire                                          [3:0] ds7_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds7_arid;
wire                                          [7:0] ds7_arlen;
wire                                                ds7_arlock;
wire                                          [2:0] ds7_arprot;
wire                                          [2:0] ds7_arsize;
wire                                                ds7_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds7_awaddr;
wire                                          [1:0] ds7_awburst;
wire                                          [3:0] ds7_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds7_awid;
wire                                          [7:0] ds7_awlen;
wire                                                ds7_awlock;
wire                                          [2:0] ds7_awprot;
wire                                          [2:0] ds7_awsize;
wire                                                ds7_awvalid;
wire                                                ds7_bready;
wire                                                ds7_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds7_wdata;
wire                                                ds7_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds7_wstrb;
wire                                                ds7_wvalid;
`endif // ATCBMC300_SLV7_SUPPORT
`ifdef ATCBMC300_SLV8_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds8_wid;
wire                                                ds8_arready;
wire                                                ds8_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds8_bid;
wire                                          [1:0] ds8_bresp;
wire                                                ds8_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds8_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds8_rid;
wire                                                ds8_rlast;
wire                                          [1:0] ds8_rresp;
wire                                                ds8_rvalid;
wire                                                ds8_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds8_araddr;
wire                                          [1:0] ds8_arburst;
wire                                          [3:0] ds8_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds8_arid;
wire                                          [7:0] ds8_arlen;
wire                                                ds8_arlock;
wire                                          [2:0] ds8_arprot;
wire                                          [2:0] ds8_arsize;
wire                                                ds8_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds8_awaddr;
wire                                          [1:0] ds8_awburst;
wire                                          [3:0] ds8_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds8_awid;
wire                                          [7:0] ds8_awlen;
wire                                                ds8_awlock;
wire                                          [2:0] ds8_awprot;
wire                                          [2:0] ds8_awsize;
wire                                                ds8_awvalid;
wire                                                ds8_bready;
wire                                                ds8_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds8_wdata;
wire                                                ds8_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds8_wstrb;
wire                                                ds8_wvalid;
`endif // ATCBMC300_SLV8_SUPPORT
`ifdef ATCBMC300_SLV9_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds9_wid;
wire                                                ds9_arready;
wire                                                ds9_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds9_bid;
wire                                          [1:0] ds9_bresp;
wire                                                ds9_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds9_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds9_rid;
wire                                                ds9_rlast;
wire                                          [1:0] ds9_rresp;
wire                                                ds9_rvalid;
wire                                                ds9_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds9_araddr;
wire                                          [1:0] ds9_arburst;
wire                                          [3:0] ds9_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds9_arid;
wire                                          [7:0] ds9_arlen;
wire                                                ds9_arlock;
wire                                          [2:0] ds9_arprot;
wire                                          [2:0] ds9_arsize;
wire                                                ds9_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds9_awaddr;
wire                                          [1:0] ds9_awburst;
wire                                          [3:0] ds9_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds9_awid;
wire                                          [7:0] ds9_awlen;
wire                                                ds9_awlock;
wire                                          [2:0] ds9_awprot;
wire                                          [2:0] ds9_awsize;
wire                                                ds9_awvalid;
wire                                                ds9_bready;
wire                                                ds9_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds9_wdata;
wire                                                ds9_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds9_wstrb;
wire                                                ds9_wvalid;
`endif // ATCBMC300_SLV9_SUPPORT
`ifdef ATCBMC300_SLV10_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds10_wid;
wire                                                ds10_arready;
wire                                                ds10_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds10_bid;
wire                                          [1:0] ds10_bresp;
wire                                                ds10_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds10_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds10_rid;
wire                                                ds10_rlast;
wire                                          [1:0] ds10_rresp;
wire                                                ds10_rvalid;
wire                                                ds10_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds10_araddr;
wire                                          [1:0] ds10_arburst;
wire                                          [3:0] ds10_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds10_arid;
wire                                          [7:0] ds10_arlen;
wire                                                ds10_arlock;
wire                                          [2:0] ds10_arprot;
wire                                          [2:0] ds10_arsize;
wire                                                ds10_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds10_awaddr;
wire                                          [1:0] ds10_awburst;
wire                                          [3:0] ds10_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds10_awid;
wire                                          [7:0] ds10_awlen;
wire                                                ds10_awlock;
wire                                          [2:0] ds10_awprot;
wire                                          [2:0] ds10_awsize;
wire                                                ds10_awvalid;
wire                                                ds10_bready;
wire                                                ds10_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds10_wdata;
wire                                                ds10_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds10_wstrb;
wire                                                ds10_wvalid;
`endif // ATCBMC300_SLV10_SUPPORT
`ifdef ATCBMC300_SLV11_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds11_wid;
wire                                                ds11_arready;
wire                                                ds11_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds11_bid;
wire                                          [1:0] ds11_bresp;
wire                                                ds11_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds11_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds11_rid;
wire                                                ds11_rlast;
wire                                          [1:0] ds11_rresp;
wire                                                ds11_rvalid;
wire                                                ds11_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds11_araddr;
wire                                          [1:0] ds11_arburst;
wire                                          [3:0] ds11_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds11_arid;
wire                                          [7:0] ds11_arlen;
wire                                                ds11_arlock;
wire                                          [2:0] ds11_arprot;
wire                                          [2:0] ds11_arsize;
wire                                                ds11_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds11_awaddr;
wire                                          [1:0] ds11_awburst;
wire                                          [3:0] ds11_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds11_awid;
wire                                          [7:0] ds11_awlen;
wire                                                ds11_awlock;
wire                                          [2:0] ds11_awprot;
wire                                          [2:0] ds11_awsize;
wire                                                ds11_awvalid;
wire                                                ds11_bready;
wire                                                ds11_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds11_wdata;
wire                                                ds11_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds11_wstrb;
wire                                                ds11_wvalid;
`endif // ATCBMC300_SLV11_SUPPORT
`ifdef ATCBMC300_SLV12_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds12_wid;
wire                                                ds12_arready;
wire                                                ds12_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds12_bid;
wire                                          [1:0] ds12_bresp;
wire                                                ds12_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds12_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds12_rid;
wire                                                ds12_rlast;
wire                                          [1:0] ds12_rresp;
wire                                                ds12_rvalid;
wire                                                ds12_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds12_araddr;
wire                                          [1:0] ds12_arburst;
wire                                          [3:0] ds12_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds12_arid;
wire                                          [7:0] ds12_arlen;
wire                                                ds12_arlock;
wire                                          [2:0] ds12_arprot;
wire                                          [2:0] ds12_arsize;
wire                                                ds12_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds12_awaddr;
wire                                          [1:0] ds12_awburst;
wire                                          [3:0] ds12_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds12_awid;
wire                                          [7:0] ds12_awlen;
wire                                                ds12_awlock;
wire                                          [2:0] ds12_awprot;
wire                                          [2:0] ds12_awsize;
wire                                                ds12_awvalid;
wire                                                ds12_bready;
wire                                                ds12_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds12_wdata;
wire                                                ds12_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds12_wstrb;
wire                                                ds12_wvalid;
`endif // ATCBMC300_SLV12_SUPPORT
`ifdef ATCBMC300_SLV13_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds13_wid;
wire                                                ds13_arready;
wire                                                ds13_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds13_bid;
wire                                          [1:0] ds13_bresp;
wire                                                ds13_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds13_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds13_rid;
wire                                                ds13_rlast;
wire                                          [1:0] ds13_rresp;
wire                                                ds13_rvalid;
wire                                                ds13_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds13_araddr;
wire                                          [1:0] ds13_arburst;
wire                                          [3:0] ds13_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds13_arid;
wire                                          [7:0] ds13_arlen;
wire                                                ds13_arlock;
wire                                          [2:0] ds13_arprot;
wire                                          [2:0] ds13_arsize;
wire                                                ds13_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds13_awaddr;
wire                                          [1:0] ds13_awburst;
wire                                          [3:0] ds13_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds13_awid;
wire                                          [7:0] ds13_awlen;
wire                                                ds13_awlock;
wire                                          [2:0] ds13_awprot;
wire                                          [2:0] ds13_awsize;
wire                                                ds13_awvalid;
wire                                                ds13_bready;
wire                                                ds13_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds13_wdata;
wire                                                ds13_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds13_wstrb;
wire                                                ds13_wvalid;
`endif // ATCBMC300_SLV13_SUPPORT
`ifdef ATCBMC300_SLV14_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds14_wid;
wire                                                ds14_arready;
wire                                                ds14_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds14_bid;
wire                                          [1:0] ds14_bresp;
wire                                                ds14_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds14_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds14_rid;
wire                                                ds14_rlast;
wire                                          [1:0] ds14_rresp;
wire                                                ds14_rvalid;
wire                                                ds14_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds14_araddr;
wire                                          [1:0] ds14_arburst;
wire                                          [3:0] ds14_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds14_arid;
wire                                          [7:0] ds14_arlen;
wire                                                ds14_arlock;
wire                                          [2:0] ds14_arprot;
wire                                          [2:0] ds14_arsize;
wire                                                ds14_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds14_awaddr;
wire                                          [1:0] ds14_awburst;
wire                                          [3:0] ds14_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds14_awid;
wire                                          [7:0] ds14_awlen;
wire                                                ds14_awlock;
wire                                          [2:0] ds14_awprot;
wire                                          [2:0] ds14_awsize;
wire                                                ds14_awvalid;
wire                                                ds14_bready;
wire                                                ds14_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds14_wdata;
wire                                                ds14_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds14_wstrb;
wire                                                ds14_wvalid;
`endif // ATCBMC300_SLV14_SUPPORT
`ifdef ATCBMC300_SLV15_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds15_wid;
wire                                                ds15_arready;
wire                                                ds15_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds15_bid;
wire                                          [1:0] ds15_bresp;
wire                                                ds15_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds15_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds15_rid;
wire                                                ds15_rlast;
wire                                          [1:0] ds15_rresp;
wire                                                ds15_rvalid;
wire                                                ds15_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds15_araddr;
wire                                          [1:0] ds15_arburst;
wire                                          [3:0] ds15_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds15_arid;
wire                                          [7:0] ds15_arlen;
wire                                                ds15_arlock;
wire                                          [2:0] ds15_arprot;
wire                                          [2:0] ds15_arsize;
wire                                                ds15_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds15_awaddr;
wire                                          [1:0] ds15_awburst;
wire                                          [3:0] ds15_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds15_awid;
wire                                          [7:0] ds15_awlen;
wire                                                ds15_awlock;
wire                                          [2:0] ds15_awprot;
wire                                          [2:0] ds15_awsize;
wire                                                ds15_awvalid;
wire                                                ds15_bready;
wire                                                ds15_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds15_wdata;
wire                                                ds15_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds15_wstrb;
wire                                                ds15_wvalid;
`endif // ATCBMC300_SLV15_SUPPORT
`ifdef ATCBMC300_SLV16_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds16_wid;
wire                                                ds16_arready;
wire                                                ds16_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds16_bid;
wire                                          [1:0] ds16_bresp;
wire                                                ds16_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds16_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds16_rid;
wire                                                ds16_rlast;
wire                                          [1:0] ds16_rresp;
wire                                                ds16_rvalid;
wire                                                ds16_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds16_araddr;
wire                                          [1:0] ds16_arburst;
wire                                          [3:0] ds16_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds16_arid;
wire                                          [7:0] ds16_arlen;
wire                                                ds16_arlock;
wire                                          [2:0] ds16_arprot;
wire                                          [2:0] ds16_arsize;
wire                                                ds16_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds16_awaddr;
wire                                          [1:0] ds16_awburst;
wire                                          [3:0] ds16_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds16_awid;
wire                                          [7:0] ds16_awlen;
wire                                                ds16_awlock;
wire                                          [2:0] ds16_awprot;
wire                                          [2:0] ds16_awsize;
wire                                                ds16_awvalid;
wire                                                ds16_bready;
wire                                                ds16_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds16_wdata;
wire                                                ds16_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds16_wstrb;
wire                                                ds16_wvalid;
`endif // ATCBMC300_SLV16_SUPPORT
`ifdef ATCBMC300_SLV17_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds17_wid;
wire                                                ds17_arready;
wire                                                ds17_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds17_bid;
wire                                          [1:0] ds17_bresp;
wire                                                ds17_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds17_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds17_rid;
wire                                                ds17_rlast;
wire                                          [1:0] ds17_rresp;
wire                                                ds17_rvalid;
wire                                                ds17_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds17_araddr;
wire                                          [1:0] ds17_arburst;
wire                                          [3:0] ds17_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds17_arid;
wire                                          [7:0] ds17_arlen;
wire                                                ds17_arlock;
wire                                          [2:0] ds17_arprot;
wire                                          [2:0] ds17_arsize;
wire                                                ds17_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds17_awaddr;
wire                                          [1:0] ds17_awburst;
wire                                          [3:0] ds17_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds17_awid;
wire                                          [7:0] ds17_awlen;
wire                                                ds17_awlock;
wire                                          [2:0] ds17_awprot;
wire                                          [2:0] ds17_awsize;
wire                                                ds17_awvalid;
wire                                                ds17_bready;
wire                                                ds17_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds17_wdata;
wire                                                ds17_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds17_wstrb;
wire                                                ds17_wvalid;
`endif // ATCBMC300_SLV17_SUPPORT
`ifdef ATCBMC300_SLV18_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds18_wid;
wire                                                ds18_arready;
wire                                                ds18_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds18_bid;
wire                                          [1:0] ds18_bresp;
wire                                                ds18_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds18_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds18_rid;
wire                                                ds18_rlast;
wire                                          [1:0] ds18_rresp;
wire                                                ds18_rvalid;
wire                                                ds18_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds18_araddr;
wire                                          [1:0] ds18_arburst;
wire                                          [3:0] ds18_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds18_arid;
wire                                          [7:0] ds18_arlen;
wire                                                ds18_arlock;
wire                                          [2:0] ds18_arprot;
wire                                          [2:0] ds18_arsize;
wire                                                ds18_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds18_awaddr;
wire                                          [1:0] ds18_awburst;
wire                                          [3:0] ds18_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds18_awid;
wire                                          [7:0] ds18_awlen;
wire                                                ds18_awlock;
wire                                          [2:0] ds18_awprot;
wire                                          [2:0] ds18_awsize;
wire                                                ds18_awvalid;
wire                                                ds18_bready;
wire                                                ds18_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds18_wdata;
wire                                                ds18_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds18_wstrb;
wire                                                ds18_wvalid;
`endif // ATCBMC300_SLV18_SUPPORT
`ifdef ATCBMC300_SLV19_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds19_wid;
wire                                                ds19_arready;
wire                                                ds19_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds19_bid;
wire                                          [1:0] ds19_bresp;
wire                                                ds19_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds19_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds19_rid;
wire                                                ds19_rlast;
wire                                          [1:0] ds19_rresp;
wire                                                ds19_rvalid;
wire                                                ds19_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds19_araddr;
wire                                          [1:0] ds19_arburst;
wire                                          [3:0] ds19_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds19_arid;
wire                                          [7:0] ds19_arlen;
wire                                                ds19_arlock;
wire                                          [2:0] ds19_arprot;
wire                                          [2:0] ds19_arsize;
wire                                                ds19_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds19_awaddr;
wire                                          [1:0] ds19_awburst;
wire                                          [3:0] ds19_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds19_awid;
wire                                          [7:0] ds19_awlen;
wire                                                ds19_awlock;
wire                                          [2:0] ds19_awprot;
wire                                          [2:0] ds19_awsize;
wire                                                ds19_awvalid;
wire                                                ds19_bready;
wire                                                ds19_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds19_wdata;
wire                                                ds19_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds19_wstrb;
wire                                                ds19_wvalid;
`endif // ATCBMC300_SLV19_SUPPORT
`ifdef ATCBMC300_SLV20_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds20_wid;
wire                                                ds20_arready;
wire                                                ds20_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds20_bid;
wire                                          [1:0] ds20_bresp;
wire                                                ds20_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds20_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds20_rid;
wire                                                ds20_rlast;
wire                                          [1:0] ds20_rresp;
wire                                                ds20_rvalid;
wire                                                ds20_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds20_araddr;
wire                                          [1:0] ds20_arburst;
wire                                          [3:0] ds20_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds20_arid;
wire                                          [7:0] ds20_arlen;
wire                                                ds20_arlock;
wire                                          [2:0] ds20_arprot;
wire                                          [2:0] ds20_arsize;
wire                                                ds20_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds20_awaddr;
wire                                          [1:0] ds20_awburst;
wire                                          [3:0] ds20_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds20_awid;
wire                                          [7:0] ds20_awlen;
wire                                                ds20_awlock;
wire                                          [2:0] ds20_awprot;
wire                                          [2:0] ds20_awsize;
wire                                                ds20_awvalid;
wire                                                ds20_bready;
wire                                                ds20_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds20_wdata;
wire                                                ds20_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds20_wstrb;
wire                                                ds20_wvalid;
`endif // ATCBMC300_SLV20_SUPPORT
`ifdef ATCBMC300_SLV21_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds21_wid;
wire                                                ds21_arready;
wire                                                ds21_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds21_bid;
wire                                          [1:0] ds21_bresp;
wire                                                ds21_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds21_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds21_rid;
wire                                                ds21_rlast;
wire                                          [1:0] ds21_rresp;
wire                                                ds21_rvalid;
wire                                                ds21_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds21_araddr;
wire                                          [1:0] ds21_arburst;
wire                                          [3:0] ds21_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds21_arid;
wire                                          [7:0] ds21_arlen;
wire                                                ds21_arlock;
wire                                          [2:0] ds21_arprot;
wire                                          [2:0] ds21_arsize;
wire                                                ds21_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds21_awaddr;
wire                                          [1:0] ds21_awburst;
wire                                          [3:0] ds21_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds21_awid;
wire                                          [7:0] ds21_awlen;
wire                                                ds21_awlock;
wire                                          [2:0] ds21_awprot;
wire                                          [2:0] ds21_awsize;
wire                                                ds21_awvalid;
wire                                                ds21_bready;
wire                                                ds21_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds21_wdata;
wire                                                ds21_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds21_wstrb;
wire                                                ds21_wvalid;
`endif // ATCBMC300_SLV21_SUPPORT
`ifdef ATCBMC300_SLV22_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds22_wid;
wire                                                ds22_arready;
wire                                                ds22_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds22_bid;
wire                                          [1:0] ds22_bresp;
wire                                                ds22_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds22_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds22_rid;
wire                                                ds22_rlast;
wire                                          [1:0] ds22_rresp;
wire                                                ds22_rvalid;
wire                                                ds22_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds22_araddr;
wire                                          [1:0] ds22_arburst;
wire                                          [3:0] ds22_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds22_arid;
wire                                          [7:0] ds22_arlen;
wire                                                ds22_arlock;
wire                                          [2:0] ds22_arprot;
wire                                          [2:0] ds22_arsize;
wire                                                ds22_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds22_awaddr;
wire                                          [1:0] ds22_awburst;
wire                                          [3:0] ds22_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds22_awid;
wire                                          [7:0] ds22_awlen;
wire                                                ds22_awlock;
wire                                          [2:0] ds22_awprot;
wire                                          [2:0] ds22_awsize;
wire                                                ds22_awvalid;
wire                                                ds22_bready;
wire                                                ds22_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds22_wdata;
wire                                                ds22_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds22_wstrb;
wire                                                ds22_wvalid;
`endif // ATCBMC300_SLV22_SUPPORT
`ifdef ATCBMC300_SLV23_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds23_wid;
wire                                                ds23_arready;
wire                                                ds23_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds23_bid;
wire                                          [1:0] ds23_bresp;
wire                                                ds23_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds23_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds23_rid;
wire                                                ds23_rlast;
wire                                          [1:0] ds23_rresp;
wire                                                ds23_rvalid;
wire                                                ds23_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds23_araddr;
wire                                          [1:0] ds23_arburst;
wire                                          [3:0] ds23_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds23_arid;
wire                                          [7:0] ds23_arlen;
wire                                                ds23_arlock;
wire                                          [2:0] ds23_arprot;
wire                                          [2:0] ds23_arsize;
wire                                                ds23_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds23_awaddr;
wire                                          [1:0] ds23_awburst;
wire                                          [3:0] ds23_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds23_awid;
wire                                          [7:0] ds23_awlen;
wire                                                ds23_awlock;
wire                                          [2:0] ds23_awprot;
wire                                          [2:0] ds23_awsize;
wire                                                ds23_awvalid;
wire                                                ds23_bready;
wire                                                ds23_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds23_wdata;
wire                                                ds23_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds23_wstrb;
wire                                                ds23_wvalid;
`endif // ATCBMC300_SLV23_SUPPORT
`ifdef ATCBMC300_SLV24_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds24_wid;
wire                                                ds24_arready;
wire                                                ds24_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds24_bid;
wire                                          [1:0] ds24_bresp;
wire                                                ds24_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds24_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds24_rid;
wire                                                ds24_rlast;
wire                                          [1:0] ds24_rresp;
wire                                                ds24_rvalid;
wire                                                ds24_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds24_araddr;
wire                                          [1:0] ds24_arburst;
wire                                          [3:0] ds24_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds24_arid;
wire                                          [7:0] ds24_arlen;
wire                                                ds24_arlock;
wire                                          [2:0] ds24_arprot;
wire                                          [2:0] ds24_arsize;
wire                                                ds24_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds24_awaddr;
wire                                          [1:0] ds24_awburst;
wire                                          [3:0] ds24_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds24_awid;
wire                                          [7:0] ds24_awlen;
wire                                                ds24_awlock;
wire                                          [2:0] ds24_awprot;
wire                                          [2:0] ds24_awsize;
wire                                                ds24_awvalid;
wire                                                ds24_bready;
wire                                                ds24_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds24_wdata;
wire                                                ds24_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds24_wstrb;
wire                                                ds24_wvalid;
`endif // ATCBMC300_SLV24_SUPPORT
`ifdef ATCBMC300_SLV25_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds25_wid;
wire                                                ds25_arready;
wire                                                ds25_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds25_bid;
wire                                          [1:0] ds25_bresp;
wire                                                ds25_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds25_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds25_rid;
wire                                                ds25_rlast;
wire                                          [1:0] ds25_rresp;
wire                                                ds25_rvalid;
wire                                                ds25_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds25_araddr;
wire                                          [1:0] ds25_arburst;
wire                                          [3:0] ds25_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds25_arid;
wire                                          [7:0] ds25_arlen;
wire                                                ds25_arlock;
wire                                          [2:0] ds25_arprot;
wire                                          [2:0] ds25_arsize;
wire                                                ds25_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds25_awaddr;
wire                                          [1:0] ds25_awburst;
wire                                          [3:0] ds25_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds25_awid;
wire                                          [7:0] ds25_awlen;
wire                                                ds25_awlock;
wire                                          [2:0] ds25_awprot;
wire                                          [2:0] ds25_awsize;
wire                                                ds25_awvalid;
wire                                                ds25_bready;
wire                                                ds25_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds25_wdata;
wire                                                ds25_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds25_wstrb;
wire                                                ds25_wvalid;
`endif // ATCBMC300_SLV25_SUPPORT
`ifdef ATCBMC300_SLV26_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds26_wid;
wire                                                ds26_arready;
wire                                                ds26_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds26_bid;
wire                                          [1:0] ds26_bresp;
wire                                                ds26_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds26_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds26_rid;
wire                                                ds26_rlast;
wire                                          [1:0] ds26_rresp;
wire                                                ds26_rvalid;
wire                                                ds26_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds26_araddr;
wire                                          [1:0] ds26_arburst;
wire                                          [3:0] ds26_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds26_arid;
wire                                          [7:0] ds26_arlen;
wire                                                ds26_arlock;
wire                                          [2:0] ds26_arprot;
wire                                          [2:0] ds26_arsize;
wire                                                ds26_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds26_awaddr;
wire                                          [1:0] ds26_awburst;
wire                                          [3:0] ds26_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds26_awid;
wire                                          [7:0] ds26_awlen;
wire                                                ds26_awlock;
wire                                          [2:0] ds26_awprot;
wire                                          [2:0] ds26_awsize;
wire                                                ds26_awvalid;
wire                                                ds26_bready;
wire                                                ds26_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds26_wdata;
wire                                                ds26_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds26_wstrb;
wire                                                ds26_wvalid;
`endif // ATCBMC300_SLV26_SUPPORT
`ifdef ATCBMC300_SLV27_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds27_wid;
wire                                                ds27_arready;
wire                                                ds27_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds27_bid;
wire                                          [1:0] ds27_bresp;
wire                                                ds27_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds27_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds27_rid;
wire                                                ds27_rlast;
wire                                          [1:0] ds27_rresp;
wire                                                ds27_rvalid;
wire                                                ds27_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds27_araddr;
wire                                          [1:0] ds27_arburst;
wire                                          [3:0] ds27_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds27_arid;
wire                                          [7:0] ds27_arlen;
wire                                                ds27_arlock;
wire                                          [2:0] ds27_arprot;
wire                                          [2:0] ds27_arsize;
wire                                                ds27_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds27_awaddr;
wire                                          [1:0] ds27_awburst;
wire                                          [3:0] ds27_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds27_awid;
wire                                          [7:0] ds27_awlen;
wire                                                ds27_awlock;
wire                                          [2:0] ds27_awprot;
wire                                          [2:0] ds27_awsize;
wire                                                ds27_awvalid;
wire                                                ds27_bready;
wire                                                ds27_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds27_wdata;
wire                                                ds27_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds27_wstrb;
wire                                                ds27_wvalid;
`endif // ATCBMC300_SLV27_SUPPORT
`ifdef ATCBMC300_SLV28_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds28_wid;
wire                                                ds28_arready;
wire                                                ds28_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds28_bid;
wire                                          [1:0] ds28_bresp;
wire                                                ds28_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds28_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds28_rid;
wire                                                ds28_rlast;
wire                                          [1:0] ds28_rresp;
wire                                                ds28_rvalid;
wire                                                ds28_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds28_araddr;
wire                                          [1:0] ds28_arburst;
wire                                          [3:0] ds28_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds28_arid;
wire                                          [7:0] ds28_arlen;
wire                                                ds28_arlock;
wire                                          [2:0] ds28_arprot;
wire                                          [2:0] ds28_arsize;
wire                                                ds28_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds28_awaddr;
wire                                          [1:0] ds28_awburst;
wire                                          [3:0] ds28_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds28_awid;
wire                                          [7:0] ds28_awlen;
wire                                                ds28_awlock;
wire                                          [2:0] ds28_awprot;
wire                                          [2:0] ds28_awsize;
wire                                                ds28_awvalid;
wire                                                ds28_bready;
wire                                                ds28_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds28_wdata;
wire                                                ds28_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds28_wstrb;
wire                                                ds28_wvalid;
`endif // ATCBMC300_SLV28_SUPPORT
`ifdef ATCBMC300_SLV29_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds29_wid;
wire                                                ds29_arready;
wire                                                ds29_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds29_bid;
wire                                          [1:0] ds29_bresp;
wire                                                ds29_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds29_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds29_rid;
wire                                                ds29_rlast;
wire                                          [1:0] ds29_rresp;
wire                                                ds29_rvalid;
wire                                                ds29_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds29_araddr;
wire                                          [1:0] ds29_arburst;
wire                                          [3:0] ds29_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds29_arid;
wire                                          [7:0] ds29_arlen;
wire                                                ds29_arlock;
wire                                          [2:0] ds29_arprot;
wire                                          [2:0] ds29_arsize;
wire                                                ds29_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds29_awaddr;
wire                                          [1:0] ds29_awburst;
wire                                          [3:0] ds29_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds29_awid;
wire                                          [7:0] ds29_awlen;
wire                                                ds29_awlock;
wire                                          [2:0] ds29_awprot;
wire                                          [2:0] ds29_awsize;
wire                                                ds29_awvalid;
wire                                                ds29_bready;
wire                                                ds29_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds29_wdata;
wire                                                ds29_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds29_wstrb;
wire                                                ds29_wvalid;
`endif // ATCBMC300_SLV29_SUPPORT
`ifdef ATCBMC300_SLV30_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds30_wid;
wire                                                ds30_arready;
wire                                                ds30_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds30_bid;
wire                                          [1:0] ds30_bresp;
wire                                                ds30_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds30_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds30_rid;
wire                                                ds30_rlast;
wire                                          [1:0] ds30_rresp;
wire                                                ds30_rvalid;
wire                                                ds30_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds30_araddr;
wire                                          [1:0] ds30_arburst;
wire                                          [3:0] ds30_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds30_arid;
wire                                          [7:0] ds30_arlen;
wire                                                ds30_arlock;
wire                                          [2:0] ds30_arprot;
wire                                          [2:0] ds30_arsize;
wire                                                ds30_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds30_awaddr;
wire                                          [1:0] ds30_awburst;
wire                                          [3:0] ds30_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds30_awid;
wire                                          [7:0] ds30_awlen;
wire                                                ds30_awlock;
wire                                          [2:0] ds30_awprot;
wire                                          [2:0] ds30_awsize;
wire                                                ds30_awvalid;
wire                                                ds30_bready;
wire                                                ds30_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds30_wdata;
wire                                                ds30_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds30_wstrb;
wire                                                ds30_wvalid;
`endif // ATCBMC300_SLV30_SUPPORT
`ifdef ATCBMC300_SLV31_SUPPORT
supply0                           [DS_ID_WIDTH-1:0] ds31_wid;
wire                                                ds31_arready;
wire                                                ds31_awready;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds31_bid;
wire                                          [1:0] ds31_bresp;
wire                                                ds31_bvalid;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds31_rdata;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds31_rid;
wire                                                ds31_rlast;
wire                                          [1:0] ds31_rresp;
wire                                                ds31_rvalid;
wire                                                ds31_wready;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds31_araddr;
wire                                          [1:0] ds31_arburst;
wire                                          [3:0] ds31_arcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds31_arid;
wire                                          [7:0] ds31_arlen;
wire                                                ds31_arlock;
wire                                          [2:0] ds31_arprot;
wire                                          [2:0] ds31_arsize;
wire                                                ds31_arvalid;
wire                  [(`ATCBMC300_ADDR_WIDTH-1):0] ds31_awaddr;
wire                                          [1:0] ds31_awburst;
wire                                          [3:0] ds31_awcache;
wire                  [(`ATCBMC300_ID_WIDTH-1)+4:0] ds31_awid;
wire                                          [7:0] ds31_awlen;
wire                                                ds31_awlock;
wire                                          [2:0] ds31_awprot;
wire                                          [2:0] ds31_awsize;
wire                                                ds31_awvalid;
wire                                                ds31_bready;
wire                                                ds31_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] ds31_wdata;
wire                                                ds31_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] ds31_wstrb;
wire                                                ds31_wvalid;
`endif // ATCBMC300_SLV31_SUPPORT
`ifdef ATCBMC300_MST1_SUPPORT
wire                               [ADDR_WIDTH-1:0] us1_araddr;
wire                                          [1:0] us1_arburst;
wire                                          [3:0] us1_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us1_arid;
wire                                          [7:0] us1_arlen;
wire                                                us1_arlock;
wire                                                us1_arlock_b1;
wire                                          [2:0] us1_arprot;
wire                                          [2:0] us1_arsize;
wire                                                us1_arvalid;
wire                               [ADDR_WIDTH-1:0] us1_awaddr;
wire                                          [1:0] us1_awburst;
wire                                          [3:0] us1_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us1_awid;
wire                                          [7:0] us1_awlen;
wire                                                us1_awlock;
wire                                                us1_awlock_b1;
wire                                          [2:0] us1_awprot;
wire                                          [2:0] us1_awsize;
wire                                                us1_awvalid;
wire                                                us1_bready;
wire                                                us1_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us1_wdata;
wire                              [US_ID_WIDTH-1:0] us1_wid;
wire                                                us1_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us1_wstrb;
wire                                                us1_wvalid;
wire                                                us1_arready;
wire                                                us1_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us1_bid;
wire                                          [1:0] us1_bresp;
wire                                                us1_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us1_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us1_rid;
wire                                                us1_rlast;
wire                                          [1:0] us1_rresp;
wire                                                us1_rvalid;
wire                                                us1_wready;
`endif // ATCBMC300_MST1_SUPPORT
`ifdef ATCBMC300_MST2_SUPPORT
wire                               [ADDR_WIDTH-1:0] us2_araddr;
wire                                          [1:0] us2_arburst;
wire                                          [3:0] us2_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us2_arid;
wire                                          [7:0] us2_arlen;
wire                                                us2_arlock;
wire                                                us2_arlock_b1;
wire                                          [2:0] us2_arprot;
wire                                          [2:0] us2_arsize;
wire                                                us2_arvalid;
wire                               [ADDR_WIDTH-1:0] us2_awaddr;
wire                                          [1:0] us2_awburst;
wire                                          [3:0] us2_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us2_awid;
wire                                          [7:0] us2_awlen;
wire                                                us2_awlock;
wire                                                us2_awlock_b1;
wire                                          [2:0] us2_awprot;
wire                                          [2:0] us2_awsize;
wire                                                us2_awvalid;
wire                                                us2_bready;
wire                                                us2_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us2_wdata;
wire                              [US_ID_WIDTH-1:0] us2_wid;
wire                                                us2_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us2_wstrb;
wire                                                us2_wvalid;
wire                                                us2_arready;
wire                                                us2_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us2_bid;
wire                                          [1:0] us2_bresp;
wire                                                us2_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us2_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us2_rid;
wire                                                us2_rlast;
wire                                          [1:0] us2_rresp;
wire                                                us2_rvalid;
wire                                                us2_wready;
`endif // ATCBMC300_MST2_SUPPORT
`ifdef ATCBMC300_MST3_SUPPORT
wire                               [ADDR_WIDTH-1:0] us3_araddr;
wire                                          [1:0] us3_arburst;
wire                                          [3:0] us3_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us3_arid;
wire                                          [7:0] us3_arlen;
wire                                                us3_arlock;
wire                                                us3_arlock_b1;
wire                                          [2:0] us3_arprot;
wire                                          [2:0] us3_arsize;
wire                                                us3_arvalid;
wire                               [ADDR_WIDTH-1:0] us3_awaddr;
wire                                          [1:0] us3_awburst;
wire                                          [3:0] us3_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us3_awid;
wire                                          [7:0] us3_awlen;
wire                                                us3_awlock;
wire                                                us3_awlock_b1;
wire                                          [2:0] us3_awprot;
wire                                          [2:0] us3_awsize;
wire                                                us3_awvalid;
wire                                                us3_bready;
wire                                                us3_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us3_wdata;
wire                              [US_ID_WIDTH-1:0] us3_wid;
wire                                                us3_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us3_wstrb;
wire                                                us3_wvalid;
wire                                                us3_arready;
wire                                                us3_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us3_bid;
wire                                          [1:0] us3_bresp;
wire                                                us3_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us3_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us3_rid;
wire                                                us3_rlast;
wire                                          [1:0] us3_rresp;
wire                                                us3_rvalid;
wire                                                us3_wready;
`endif // ATCBMC300_MST3_SUPPORT
`ifdef ATCBMC300_MST4_SUPPORT
wire                               [ADDR_WIDTH-1:0] us4_araddr;
wire                                          [1:0] us4_arburst;
wire                                          [3:0] us4_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us4_arid;
wire                                          [7:0] us4_arlen;
wire                                                us4_arlock;
wire                                                us4_arlock_b1;
wire                                          [2:0] us4_arprot;
wire                                          [2:0] us4_arsize;
wire                                                us4_arvalid;
wire                               [ADDR_WIDTH-1:0] us4_awaddr;
wire                                          [1:0] us4_awburst;
wire                                          [3:0] us4_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us4_awid;
wire                                          [7:0] us4_awlen;
wire                                                us4_awlock;
wire                                                us4_awlock_b1;
wire                                          [2:0] us4_awprot;
wire                                          [2:0] us4_awsize;
wire                                                us4_awvalid;
wire                                                us4_bready;
wire                                                us4_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us4_wdata;
wire                              [US_ID_WIDTH-1:0] us4_wid;
wire                                                us4_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us4_wstrb;
wire                                                us4_wvalid;
wire                                                us4_arready;
wire                                                us4_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us4_bid;
wire                                          [1:0] us4_bresp;
wire                                                us4_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us4_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us4_rid;
wire                                                us4_rlast;
wire                                          [1:0] us4_rresp;
wire                                                us4_rvalid;
wire                                                us4_wready;
`endif // ATCBMC300_MST4_SUPPORT
`ifdef ATCBMC300_MST5_SUPPORT
wire                               [ADDR_WIDTH-1:0] us5_araddr;
wire                                          [1:0] us5_arburst;
wire                                          [3:0] us5_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us5_arid;
wire                                          [7:0] us5_arlen;
wire                                                us5_arlock;
wire                                                us5_arlock_b1;
wire                                          [2:0] us5_arprot;
wire                                          [2:0] us5_arsize;
wire                                                us5_arvalid;
wire                               [ADDR_WIDTH-1:0] us5_awaddr;
wire                                          [1:0] us5_awburst;
wire                                          [3:0] us5_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us5_awid;
wire                                          [7:0] us5_awlen;
wire                                                us5_awlock;
wire                                                us5_awlock_b1;
wire                                          [2:0] us5_awprot;
wire                                          [2:0] us5_awsize;
wire                                                us5_awvalid;
wire                                                us5_bready;
wire                                                us5_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us5_wdata;
wire                              [US_ID_WIDTH-1:0] us5_wid;
wire                                                us5_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us5_wstrb;
wire                                                us5_wvalid;
wire                                                us5_arready;
wire                                                us5_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us5_bid;
wire                                          [1:0] us5_bresp;
wire                                                us5_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us5_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us5_rid;
wire                                                us5_rlast;
wire                                          [1:0] us5_rresp;
wire                                                us5_rvalid;
wire                                                us5_wready;
`endif // ATCBMC300_MST5_SUPPORT
`ifdef ATCBMC300_MST6_SUPPORT
wire                               [ADDR_WIDTH-1:0] us6_araddr;
wire                                          [1:0] us6_arburst;
wire                                          [3:0] us6_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us6_arid;
wire                                          [7:0] us6_arlen;
wire                                                us6_arlock;
wire                                                us6_arlock_b1;
wire                                          [2:0] us6_arprot;
wire                                          [2:0] us6_arsize;
wire                                                us6_arvalid;
wire                               [ADDR_WIDTH-1:0] us6_awaddr;
wire                                          [1:0] us6_awburst;
wire                                          [3:0] us6_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us6_awid;
wire                                          [7:0] us6_awlen;
wire                                                us6_awlock;
wire                                                us6_awlock_b1;
wire                                          [2:0] us6_awprot;
wire                                          [2:0] us6_awsize;
wire                                                us6_awvalid;
wire                                                us6_bready;
wire                                                us6_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us6_wdata;
wire                              [US_ID_WIDTH-1:0] us6_wid;
wire                                                us6_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us6_wstrb;
wire                                                us6_wvalid;
wire                                                us6_arready;
wire                                                us6_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us6_bid;
wire                                          [1:0] us6_bresp;
wire                                                us6_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us6_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us6_rid;
wire                                                us6_rlast;
wire                                          [1:0] us6_rresp;
wire                                                us6_rvalid;
wire                                                us6_wready;
`endif // ATCBMC300_MST6_SUPPORT
`ifdef ATCBMC300_MST7_SUPPORT
wire                               [ADDR_WIDTH-1:0] us7_araddr;
wire                                          [1:0] us7_arburst;
wire                                          [3:0] us7_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us7_arid;
wire                                          [7:0] us7_arlen;
wire                                                us7_arlock;
wire                                                us7_arlock_b1;
wire                                          [2:0] us7_arprot;
wire                                          [2:0] us7_arsize;
wire                                                us7_arvalid;
wire                               [ADDR_WIDTH-1:0] us7_awaddr;
wire                                          [1:0] us7_awburst;
wire                                          [3:0] us7_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us7_awid;
wire                                          [7:0] us7_awlen;
wire                                                us7_awlock;
wire                                                us7_awlock_b1;
wire                                          [2:0] us7_awprot;
wire                                          [2:0] us7_awsize;
wire                                                us7_awvalid;
wire                                                us7_bready;
wire                                                us7_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us7_wdata;
wire                              [US_ID_WIDTH-1:0] us7_wid;
wire                                                us7_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us7_wstrb;
wire                                                us7_wvalid;
wire                                                us7_arready;
wire                                                us7_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us7_bid;
wire                                          [1:0] us7_bresp;
wire                                                us7_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us7_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us7_rid;
wire                                                us7_rlast;
wire                                          [1:0] us7_rresp;
wire                                                us7_rvalid;
wire                                                us7_wready;
`endif // ATCBMC300_MST7_SUPPORT
`ifdef ATCBMC300_MST8_SUPPORT
wire                               [ADDR_WIDTH-1:0] us8_araddr;
wire                                          [1:0] us8_arburst;
wire                                          [3:0] us8_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us8_arid;
wire                                          [7:0] us8_arlen;
wire                                                us8_arlock;
wire                                                us8_arlock_b1;
wire                                          [2:0] us8_arprot;
wire                                          [2:0] us8_arsize;
wire                                                us8_arvalid;
wire                               [ADDR_WIDTH-1:0] us8_awaddr;
wire                                          [1:0] us8_awburst;
wire                                          [3:0] us8_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us8_awid;
wire                                          [7:0] us8_awlen;
wire                                                us8_awlock;
wire                                                us8_awlock_b1;
wire                                          [2:0] us8_awprot;
wire                                          [2:0] us8_awsize;
wire                                                us8_awvalid;
wire                                                us8_bready;
wire                                                us8_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us8_wdata;
wire                              [US_ID_WIDTH-1:0] us8_wid;
wire                                                us8_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us8_wstrb;
wire                                                us8_wvalid;
wire                                                us8_arready;
wire                                                us8_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us8_bid;
wire                                          [1:0] us8_bresp;
wire                                                us8_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us8_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us8_rid;
wire                                                us8_rlast;
wire                                          [1:0] us8_rresp;
wire                                                us8_rvalid;
wire                                                us8_wready;
`endif // ATCBMC300_MST8_SUPPORT
`ifdef ATCBMC300_MST9_SUPPORT
wire                               [ADDR_WIDTH-1:0] us9_araddr;
wire                                          [1:0] us9_arburst;
wire                                          [3:0] us9_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us9_arid;
wire                                          [7:0] us9_arlen;
wire                                                us9_arlock;
wire                                                us9_arlock_b1;
wire                                          [2:0] us9_arprot;
wire                                          [2:0] us9_arsize;
wire                                                us9_arvalid;
wire                               [ADDR_WIDTH-1:0] us9_awaddr;
wire                                          [1:0] us9_awburst;
wire                                          [3:0] us9_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us9_awid;
wire                                          [7:0] us9_awlen;
wire                                                us9_awlock;
wire                                                us9_awlock_b1;
wire                                          [2:0] us9_awprot;
wire                                          [2:0] us9_awsize;
wire                                                us9_awvalid;
wire                                                us9_bready;
wire                                                us9_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us9_wdata;
wire                              [US_ID_WIDTH-1:0] us9_wid;
wire                                                us9_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us9_wstrb;
wire                                                us9_wvalid;
wire                                                us9_arready;
wire                                                us9_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us9_bid;
wire                                          [1:0] us9_bresp;
wire                                                us9_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us9_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us9_rid;
wire                                                us9_rlast;
wire                                          [1:0] us9_rresp;
wire                                                us9_rvalid;
wire                                                us9_wready;
`endif // ATCBMC300_MST9_SUPPORT
`ifdef ATCBMC300_MST10_SUPPORT
wire                               [ADDR_WIDTH-1:0] us10_araddr;
wire                                          [1:0] us10_arburst;
wire                                          [3:0] us10_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us10_arid;
wire                                          [7:0] us10_arlen;
wire                                                us10_arlock;
wire                                                us10_arlock_b1;
wire                                          [2:0] us10_arprot;
wire                                          [2:0] us10_arsize;
wire                                                us10_arvalid;
wire                               [ADDR_WIDTH-1:0] us10_awaddr;
wire                                          [1:0] us10_awburst;
wire                                          [3:0] us10_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us10_awid;
wire                                          [7:0] us10_awlen;
wire                                                us10_awlock;
wire                                                us10_awlock_b1;
wire                                          [2:0] us10_awprot;
wire                                          [2:0] us10_awsize;
wire                                                us10_awvalid;
wire                                                us10_bready;
wire                                                us10_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us10_wdata;
wire                              [US_ID_WIDTH-1:0] us10_wid;
wire                                                us10_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us10_wstrb;
wire                                                us10_wvalid;
wire                                                us10_arready;
wire                                                us10_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us10_bid;
wire                                          [1:0] us10_bresp;
wire                                                us10_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us10_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us10_rid;
wire                                                us10_rlast;
wire                                          [1:0] us10_rresp;
wire                                                us10_rvalid;
wire                                                us10_wready;
`endif // ATCBMC300_MST10_SUPPORT
`ifdef ATCBMC300_MST11_SUPPORT
wire                               [ADDR_WIDTH-1:0] us11_araddr;
wire                                          [1:0] us11_arburst;
wire                                          [3:0] us11_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us11_arid;
wire                                          [7:0] us11_arlen;
wire                                                us11_arlock;
wire                                                us11_arlock_b1;
wire                                          [2:0] us11_arprot;
wire                                          [2:0] us11_arsize;
wire                                                us11_arvalid;
wire                               [ADDR_WIDTH-1:0] us11_awaddr;
wire                                          [1:0] us11_awburst;
wire                                          [3:0] us11_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us11_awid;
wire                                          [7:0] us11_awlen;
wire                                                us11_awlock;
wire                                                us11_awlock_b1;
wire                                          [2:0] us11_awprot;
wire                                          [2:0] us11_awsize;
wire                                                us11_awvalid;
wire                                                us11_bready;
wire                                                us11_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us11_wdata;
wire                              [US_ID_WIDTH-1:0] us11_wid;
wire                                                us11_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us11_wstrb;
wire                                                us11_wvalid;
wire                                                us11_arready;
wire                                                us11_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us11_bid;
wire                                          [1:0] us11_bresp;
wire                                                us11_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us11_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us11_rid;
wire                                                us11_rlast;
wire                                          [1:0] us11_rresp;
wire                                                us11_rvalid;
wire                                                us11_wready;
`endif // ATCBMC300_MST11_SUPPORT
`ifdef ATCBMC300_MST12_SUPPORT
wire                               [ADDR_WIDTH-1:0] us12_araddr;
wire                                          [1:0] us12_arburst;
wire                                          [3:0] us12_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us12_arid;
wire                                          [7:0] us12_arlen;
wire                                                us12_arlock;
wire                                                us12_arlock_b1;
wire                                          [2:0] us12_arprot;
wire                                          [2:0] us12_arsize;
wire                                                us12_arvalid;
wire                               [ADDR_WIDTH-1:0] us12_awaddr;
wire                                          [1:0] us12_awburst;
wire                                          [3:0] us12_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us12_awid;
wire                                          [7:0] us12_awlen;
wire                                                us12_awlock;
wire                                                us12_awlock_b1;
wire                                          [2:0] us12_awprot;
wire                                          [2:0] us12_awsize;
wire                                                us12_awvalid;
wire                                                us12_bready;
wire                                                us12_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us12_wdata;
wire                              [US_ID_WIDTH-1:0] us12_wid;
wire                                                us12_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us12_wstrb;
wire                                                us12_wvalid;
wire                                                us12_arready;
wire                                                us12_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us12_bid;
wire                                          [1:0] us12_bresp;
wire                                                us12_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us12_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us12_rid;
wire                                                us12_rlast;
wire                                          [1:0] us12_rresp;
wire                                                us12_rvalid;
wire                                                us12_wready;
`endif // ATCBMC300_MST12_SUPPORT
`ifdef ATCBMC300_MST13_SUPPORT
wire                               [ADDR_WIDTH-1:0] us13_araddr;
wire                                          [1:0] us13_arburst;
wire                                          [3:0] us13_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us13_arid;
wire                                          [7:0] us13_arlen;
wire                                                us13_arlock;
wire                                                us13_arlock_b1;
wire                                          [2:0] us13_arprot;
wire                                          [2:0] us13_arsize;
wire                                                us13_arvalid;
wire                               [ADDR_WIDTH-1:0] us13_awaddr;
wire                                          [1:0] us13_awburst;
wire                                          [3:0] us13_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us13_awid;
wire                                          [7:0] us13_awlen;
wire                                                us13_awlock;
wire                                                us13_awlock_b1;
wire                                          [2:0] us13_awprot;
wire                                          [2:0] us13_awsize;
wire                                                us13_awvalid;
wire                                                us13_bready;
wire                                                us13_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us13_wdata;
wire                              [US_ID_WIDTH-1:0] us13_wid;
wire                                                us13_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us13_wstrb;
wire                                                us13_wvalid;
wire                                                us13_arready;
wire                                                us13_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us13_bid;
wire                                          [1:0] us13_bresp;
wire                                                us13_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us13_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us13_rid;
wire                                                us13_rlast;
wire                                          [1:0] us13_rresp;
wire                                                us13_rvalid;
wire                                                us13_wready;
`endif // ATCBMC300_MST13_SUPPORT
`ifdef ATCBMC300_MST14_SUPPORT
wire                               [ADDR_WIDTH-1:0] us14_araddr;
wire                                          [1:0] us14_arburst;
wire                                          [3:0] us14_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us14_arid;
wire                                          [7:0] us14_arlen;
wire                                                us14_arlock;
wire                                                us14_arlock_b1;
wire                                          [2:0] us14_arprot;
wire                                          [2:0] us14_arsize;
wire                                                us14_arvalid;
wire                               [ADDR_WIDTH-1:0] us14_awaddr;
wire                                          [1:0] us14_awburst;
wire                                          [3:0] us14_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us14_awid;
wire                                          [7:0] us14_awlen;
wire                                                us14_awlock;
wire                                                us14_awlock_b1;
wire                                          [2:0] us14_awprot;
wire                                          [2:0] us14_awsize;
wire                                                us14_awvalid;
wire                                                us14_bready;
wire                                                us14_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us14_wdata;
wire                              [US_ID_WIDTH-1:0] us14_wid;
wire                                                us14_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us14_wstrb;
wire                                                us14_wvalid;
wire                                                us14_arready;
wire                                                us14_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us14_bid;
wire                                          [1:0] us14_bresp;
wire                                                us14_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us14_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us14_rid;
wire                                                us14_rlast;
wire                                          [1:0] us14_rresp;
wire                                                us14_rvalid;
wire                                                us14_wready;
`endif // ATCBMC300_MST14_SUPPORT
`ifdef ATCBMC300_MST15_SUPPORT
wire                               [ADDR_WIDTH-1:0] us15_araddr;
wire                                          [1:0] us15_arburst;
wire                                          [3:0] us15_arcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us15_arid;
wire                                          [7:0] us15_arlen;
wire                                                us15_arlock;
wire                                                us15_arlock_b1;
wire                                          [2:0] us15_arprot;
wire                                          [2:0] us15_arsize;
wire                                                us15_arvalid;
wire                               [ADDR_WIDTH-1:0] us15_awaddr;
wire                                          [1:0] us15_awburst;
wire                                          [3:0] us15_awcache;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us15_awid;
wire                                          [7:0] us15_awlen;
wire                                                us15_awlock;
wire                                                us15_awlock_b1;
wire                                          [2:0] us15_awprot;
wire                                          [2:0] us15_awsize;
wire                                                us15_awvalid;
wire                                                us15_bready;
wire                                                us15_rready;
wire                  [(`ATCBMC300_DATA_WIDTH-1):0] us15_wdata;
wire                              [US_ID_WIDTH-1:0] us15_wid;
wire                                                us15_wlast;
wire        [(((`ATCBMC300_DATA_WIDTH-1)+1)/8)-1:0] us15_wstrb;
wire                                                us15_wvalid;
wire                                                us15_arready;
wire                                                us15_awready;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us15_bid;
wire                                          [1:0] us15_bresp;
wire                                                us15_bvalid;
wire                    [`ATCBMC300_DATA_WIDTH-1:0] us15_rdata;
wire                    [(`ATCBMC300_ID_WIDTH-1):0] us15_rid;
wire                                                us15_rlast;
wire                                          [1:0] us15_rresp;
wire                                                us15_rvalid;
wire                                                us15_wready;
`endif // ATCBMC300_MST15_SUPPORT
`ifdef NDS_AXI_AWREGION_SUPPORT
wire                                          [3:0] awregion;
`endif // NDS_AXI_AWREGION_SUPPORT
`ifdef NDS_AXI_AWQOS_SUPPORT
wire                                          [3:0] awqos;
`endif // NDS_AXI_AWQOS_SUPPORT
`ifdef NDS_AXI_AWUSER_SUPPORT
wire                                         [-1:0] awuser;
`endif // NDS_AXI_AWUSER_SUPPORT
`ifdef NDS_AXI_WUSER_SUPPORT
wire                                         [-1:0] wuser;
`endif // NDS_AXI_WUSER_SUPPORT
`ifdef NDS_AXI_BUSER_SUPPORT
wire                                         [-1:0] buser;
`endif // NDS_AXI_BUSER_SUPPORT
`ifdef NDS_AXI_ARREGION_SUPPORT
wire                                          [3:0] arregion;
`endif // NDS_AXI_ARREGION_SUPPORT
`ifdef NDS_AXI_ARQOS_SUPPORT
wire                                          [3:0] arqos;
`endif // NDS_AXI_ARQOS_SUPPORT
`ifdef NDS_AXI_ARUSER_SUPPORT
wire                                         [-1:0] aruser;
`endif // NDS_AXI_ARUSER_SUPPORT
`ifdef NDS_AXI_RUSER_SUPPORT
wire                                         [-1:0] ruser;
`endif // NDS_AXI_RUSER_SUPPORT
wire                                                aclk;
wire                                                aresetn;

`ifdef NDS_SCOREBOARD_EN
// scoreboard
blk_scb  blk_scb();

`ifdef ATCBMC300_MST0_SUPPORT
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master0.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST1_SUPPORT
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master1.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST2_SUPPORT
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master2.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST3_SUPPORT
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master3.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST4_SUPPORT
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master4.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST5_SUPPORT
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master5.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST6_SUPPORT
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master6.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST7_SUPPORT
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master7.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST8_SUPPORT
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master8.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST9_SUPPORT
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master9.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST10_SUPPORT
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master10.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST11_SUPPORT
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master11.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST12_SUPPORT
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master12.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST13_SUPPORT
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master13.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST14_SUPPORT
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master14.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif
`ifdef ATCBMC300_MST15_SUPPORT
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.ID_WIDTH = US_ID_WIDTH;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.EXCLUSIVE_TEST = 1'b0;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_master15.scb_axim_mon.CAPTURE_ID = 1'b1;
`endif

`ifdef ATCBMC300_SLV1_SUPPORT
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave1.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave1.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV2_SUPPORT
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave2.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave2.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV3_SUPPORT
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave3.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave3.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV4_SUPPORT
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave4.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave4.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV5_SUPPORT
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave5.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave5.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV6_SUPPORT
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave6.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave6.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV7_SUPPORT
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave7.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave7.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV8_SUPPORT
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave8.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave8.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV9_SUPPORT
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave9.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave9.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV10_SUPPORT
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave10.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave10.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV11_SUPPORT
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave11.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave11.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV12_SUPPORT
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave12.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave12.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV13_SUPPORT
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave13.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave13.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV14_SUPPORT
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave14.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave14.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV15_SUPPORT
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave15.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave15.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV16_SUPPORT
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave16.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave16.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV17_SUPPORT
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave17.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave17.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV18_SUPPORT
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave18.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave18.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV19_SUPPORT
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave19.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave19.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV20_SUPPORT
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave20.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave20.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV21_SUPPORT
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave21.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave21.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV22_SUPPORT
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave22.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave22.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV23_SUPPORT
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave23.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave23.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV24_SUPPORT
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave24.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave24.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV25_SUPPORT
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave25.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave25.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV26_SUPPORT
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave26.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave26.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV27_SUPPORT
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave27.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave27.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV28_SUPPORT
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave28.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave28.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV29_SUPPORT
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave29.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave29.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV30_SUPPORT
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave30.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave30.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`ifdef ATCBMC300_SLV31_SUPPORT
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.ADDR_WIDTH = ADDR_WIDTH;
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.DATA_WIDTH_SIZE = DATA_SIZE;
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.SCB_ID_WIDTH = 8;
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.ID_WIDTH = DS_ID_WIDTH;
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.AXI4 = 1'b1;
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.CAPTURE_LOCK = 1'b1;
defparam `NDS_SYSTEM.axi_slave31.scb_axis_mon.CAPTURE_ID = 1'b1;
`ifdef NDS_AXI_SLAVE_PAT	// The linter doesn't see NDS_AXI_SLAVE_PAT.
defparam `NDS_SYSTEM.axi_slave31.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
`endif
`endif
`endif // NDS_SCOREBOARD_EN


atcbmc300 bmc300 (
`ifdef ATCBMC300_MST0_SUPPORT
	.us0_araddr  (us0_araddr  ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_arburst (us0_arburst ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arcache (us0_arcache ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arid    (us0_arid    ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arlen   (us0_arlen   ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arlock  (us0_arlock  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arprot  (us0_arprot  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arready (us0_arready ), // (bmc300) => (axi_master0,axi_monitor_m0,bench)
	.us0_arsize  (us0_arsize  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_arvalid (us0_arvalid ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_awaddr  (us0_awaddr  ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_awburst (us0_awburst ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awcache (us0_awcache ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awid    (us0_awid    ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awlen   (us0_awlen   ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awlock  (us0_awlock  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awprot  (us0_awprot  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awready (us0_awready ), // (bmc300) => (axi_master0,axi_monitor_m0,bench)
	.us0_awsize  (us0_awsize  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_awvalid (us0_awvalid ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_bid     (us0_bid     ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_bready  (us0_bready  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_bresp   (us0_bresp   ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_bvalid  (us0_bvalid  ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_rdata   (us0_rdata   ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_rid     (us0_rid     ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_rlast   (us0_rlast   ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_rready  (us0_rready  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_rresp   (us0_rresp   ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_rvalid  (us0_rvalid  ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_wdata   (us0_wdata   ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_wlast   (us0_wlast   ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_wready  (us0_wready  ), // (bmc300) => (axi_master0,axi_monitor_m0)
	.us0_wstrb   (us0_wstrb   ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.us0_wvalid  (us0_wvalid  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
`endif // ATCBMC300_MST0_SUPPORT
`ifdef ATCBMC300_SLV1_SUPPORT
	.ds1_araddr  (ds1_araddr  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arburst (ds1_arburst ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arcache (ds1_arcache ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arid    (ds1_arid    ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arlen   (ds1_arlen   ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arlock  (ds1_arlock  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arprot  (ds1_arprot  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arready (ds1_arready ), // (axi_monitor_s1,bench,bmc300) <= (axi_slave1)
	.ds1_arsize  (ds1_arsize  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_arvalid (ds1_arvalid ), // (bmc300) => (axi_monitor_s1,axi_slave1,bench)
	.ds1_awaddr  (ds1_awaddr  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awburst (ds1_awburst ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awcache (ds1_awcache ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awid    (ds1_awid    ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awlen   (ds1_awlen   ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awlock  (ds1_awlock  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awprot  (ds1_awprot  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awready (ds1_awready ), // (axi_monitor_s1,bench,bmc300) <= (axi_slave1)
	.ds1_awsize  (ds1_awsize  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_awvalid (ds1_awvalid ), // (bmc300) => (axi_monitor_s1,axi_slave1,bench)
	.ds1_bid     (ds1_bid     ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_bready  (ds1_bready  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_bresp   (ds1_bresp   ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_bvalid  (ds1_bvalid  ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_rdata   (ds1_rdata   ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_rid     (ds1_rid     ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_rlast   (ds1_rlast   ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_rready  (ds1_rready  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_rresp   (ds1_rresp   ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_rvalid  (ds1_rvalid  ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_wdata   (ds1_wdata   ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_wlast   (ds1_wlast   ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_wready  (ds1_wready  ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.ds1_wstrb   (ds1_wstrb   ), // (bmc300) => (axi_monitor_s1,axi_slave1)
	.ds1_wvalid  (ds1_wvalid  ), // (bmc300) => (axi_monitor_s1,axi_slave1)
`endif // ATCBMC300_SLV1_SUPPORT
`ifdef ATCBMC300_SLV2_SUPPORT
	.ds2_araddr  (ds2_araddr  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arburst (ds2_arburst ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arcache (ds2_arcache ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arid    (ds2_arid    ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arlen   (ds2_arlen   ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arlock  (ds2_arlock  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arprot  (ds2_arprot  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arready (ds2_arready ), // (axi_monitor_s2,bench,bmc300) <= (axi_slave2)
	.ds2_arsize  (ds2_arsize  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_arvalid (ds2_arvalid ), // (bmc300) => (axi_monitor_s2,axi_slave2,bench)
	.ds2_awaddr  (ds2_awaddr  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awburst (ds2_awburst ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awcache (ds2_awcache ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awid    (ds2_awid    ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awlen   (ds2_awlen   ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awlock  (ds2_awlock  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awprot  (ds2_awprot  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awready (ds2_awready ), // (axi_monitor_s2,bench,bmc300) <= (axi_slave2)
	.ds2_awsize  (ds2_awsize  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_awvalid (ds2_awvalid ), // (bmc300) => (axi_monitor_s2,axi_slave2,bench)
	.ds2_bid     (ds2_bid     ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_bready  (ds2_bready  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_bresp   (ds2_bresp   ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_bvalid  (ds2_bvalid  ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_rdata   (ds2_rdata   ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_rid     (ds2_rid     ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_rlast   (ds2_rlast   ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_rready  (ds2_rready  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_rresp   (ds2_rresp   ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_rvalid  (ds2_rvalid  ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_wdata   (ds2_wdata   ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_wlast   (ds2_wlast   ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_wready  (ds2_wready  ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.ds2_wstrb   (ds2_wstrb   ), // (bmc300) => (axi_monitor_s2,axi_slave2)
	.ds2_wvalid  (ds2_wvalid  ), // (bmc300) => (axi_monitor_s2,axi_slave2)
`endif // ATCBMC300_SLV2_SUPPORT
`ifdef ATCBMC300_SLV3_SUPPORT
	.ds3_araddr  (ds3_araddr  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arburst (ds3_arburst ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arcache (ds3_arcache ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arid    (ds3_arid    ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arlen   (ds3_arlen   ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arlock  (ds3_arlock  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arprot  (ds3_arprot  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arready (ds3_arready ), // (axi_monitor_s3,bench,bmc300) <= (axi_slave3)
	.ds3_arsize  (ds3_arsize  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_arvalid (ds3_arvalid ), // (bmc300) => (axi_monitor_s3,axi_slave3,bench)
	.ds3_awaddr  (ds3_awaddr  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awburst (ds3_awburst ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awcache (ds3_awcache ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awid    (ds3_awid    ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awlen   (ds3_awlen   ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awlock  (ds3_awlock  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awprot  (ds3_awprot  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awready (ds3_awready ), // (axi_monitor_s3,bench,bmc300) <= (axi_slave3)
	.ds3_awsize  (ds3_awsize  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_awvalid (ds3_awvalid ), // (bmc300) => (axi_monitor_s3,axi_slave3,bench)
	.ds3_bid     (ds3_bid     ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_bready  (ds3_bready  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_bresp   (ds3_bresp   ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_bvalid  (ds3_bvalid  ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_rdata   (ds3_rdata   ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_rid     (ds3_rid     ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_rlast   (ds3_rlast   ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_rready  (ds3_rready  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_rresp   (ds3_rresp   ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_rvalid  (ds3_rvalid  ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_wdata   (ds3_wdata   ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_wlast   (ds3_wlast   ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_wready  (ds3_wready  ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.ds3_wstrb   (ds3_wstrb   ), // (bmc300) => (axi_monitor_s3,axi_slave3)
	.ds3_wvalid  (ds3_wvalid  ), // (bmc300) => (axi_monitor_s3,axi_slave3)
`endif // ATCBMC300_SLV3_SUPPORT
`ifdef ATCBMC300_SLV4_SUPPORT
	.ds4_araddr  (ds4_araddr  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arburst (ds4_arburst ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arcache (ds4_arcache ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arid    (ds4_arid    ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arlen   (ds4_arlen   ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arlock  (ds4_arlock  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arprot  (ds4_arprot  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arready (ds4_arready ), // (axi_monitor_s4,bench,bmc300) <= (axi_slave4)
	.ds4_arsize  (ds4_arsize  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_arvalid (ds4_arvalid ), // (bmc300) => (axi_monitor_s4,axi_slave4,bench)
	.ds4_awaddr  (ds4_awaddr  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awburst (ds4_awburst ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awcache (ds4_awcache ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awid    (ds4_awid    ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awlen   (ds4_awlen   ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awlock  (ds4_awlock  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awprot  (ds4_awprot  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awready (ds4_awready ), // (axi_monitor_s4,bench,bmc300) <= (axi_slave4)
	.ds4_awsize  (ds4_awsize  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_awvalid (ds4_awvalid ), // (bmc300) => (axi_monitor_s4,axi_slave4,bench)
	.ds4_bid     (ds4_bid     ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_bready  (ds4_bready  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_bresp   (ds4_bresp   ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_bvalid  (ds4_bvalid  ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_rdata   (ds4_rdata   ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_rid     (ds4_rid     ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_rlast   (ds4_rlast   ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_rready  (ds4_rready  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_rresp   (ds4_rresp   ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_rvalid  (ds4_rvalid  ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_wdata   (ds4_wdata   ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_wlast   (ds4_wlast   ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_wready  (ds4_wready  ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.ds4_wstrb   (ds4_wstrb   ), // (bmc300) => (axi_monitor_s4,axi_slave4)
	.ds4_wvalid  (ds4_wvalid  ), // (bmc300) => (axi_monitor_s4,axi_slave4)
`endif // ATCBMC300_SLV4_SUPPORT
`ifdef ATCBMC300_SLV5_SUPPORT
	.ds5_araddr  (ds5_araddr  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arburst (ds5_arburst ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arcache (ds5_arcache ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arid    (ds5_arid    ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arlen   (ds5_arlen   ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arlock  (ds5_arlock  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arprot  (ds5_arprot  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arready (ds5_arready ), // (axi_monitor_s5,bench,bmc300) <= (axi_slave5)
	.ds5_arsize  (ds5_arsize  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_arvalid (ds5_arvalid ), // (bmc300) => (axi_monitor_s5,axi_slave5,bench)
	.ds5_awaddr  (ds5_awaddr  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awburst (ds5_awburst ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awcache (ds5_awcache ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awid    (ds5_awid    ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awlen   (ds5_awlen   ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awlock  (ds5_awlock  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awprot  (ds5_awprot  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awready (ds5_awready ), // (axi_monitor_s5,bench,bmc300) <= (axi_slave5)
	.ds5_awsize  (ds5_awsize  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_awvalid (ds5_awvalid ), // (bmc300) => (axi_monitor_s5,axi_slave5,bench)
	.ds5_bid     (ds5_bid     ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_bready  (ds5_bready  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_bresp   (ds5_bresp   ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_bvalid  (ds5_bvalid  ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_rdata   (ds5_rdata   ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_rid     (ds5_rid     ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_rlast   (ds5_rlast   ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_rready  (ds5_rready  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_rresp   (ds5_rresp   ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_rvalid  (ds5_rvalid  ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_wdata   (ds5_wdata   ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_wlast   (ds5_wlast   ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_wready  (ds5_wready  ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.ds5_wstrb   (ds5_wstrb   ), // (bmc300) => (axi_monitor_s5,axi_slave5)
	.ds5_wvalid  (ds5_wvalid  ), // (bmc300) => (axi_monitor_s5,axi_slave5)
`endif // ATCBMC300_SLV5_SUPPORT
`ifdef ATCBMC300_SLV6_SUPPORT
	.ds6_araddr  (ds6_araddr  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arburst (ds6_arburst ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arcache (ds6_arcache ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arid    (ds6_arid    ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arlen   (ds6_arlen   ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arlock  (ds6_arlock  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arprot  (ds6_arprot  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arready (ds6_arready ), // (axi_monitor_s6,bench,bmc300) <= (axi_slave6)
	.ds6_arsize  (ds6_arsize  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_arvalid (ds6_arvalid ), // (bmc300) => (axi_monitor_s6,axi_slave6,bench)
	.ds6_awaddr  (ds6_awaddr  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awburst (ds6_awburst ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awcache (ds6_awcache ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awid    (ds6_awid    ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awlen   (ds6_awlen   ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awlock  (ds6_awlock  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awprot  (ds6_awprot  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awready (ds6_awready ), // (axi_monitor_s6,bench,bmc300) <= (axi_slave6)
	.ds6_awsize  (ds6_awsize  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_awvalid (ds6_awvalid ), // (bmc300) => (axi_monitor_s6,axi_slave6,bench)
	.ds6_bid     (ds6_bid     ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_bready  (ds6_bready  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_bresp   (ds6_bresp   ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_bvalid  (ds6_bvalid  ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_rdata   (ds6_rdata   ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_rid     (ds6_rid     ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_rlast   (ds6_rlast   ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_rready  (ds6_rready  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_rresp   (ds6_rresp   ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_rvalid  (ds6_rvalid  ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_wdata   (ds6_wdata   ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_wlast   (ds6_wlast   ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_wready  (ds6_wready  ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.ds6_wstrb   (ds6_wstrb   ), // (bmc300) => (axi_monitor_s6,axi_slave6)
	.ds6_wvalid  (ds6_wvalid  ), // (bmc300) => (axi_monitor_s6,axi_slave6)
`endif // ATCBMC300_SLV6_SUPPORT
`ifdef ATCBMC300_SLV7_SUPPORT
	.ds7_araddr  (ds7_araddr  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arburst (ds7_arburst ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arcache (ds7_arcache ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arid    (ds7_arid    ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arlen   (ds7_arlen   ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arlock  (ds7_arlock  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arprot  (ds7_arprot  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arready (ds7_arready ), // (axi_monitor_s7,bench,bmc300) <= (axi_slave7)
	.ds7_arsize  (ds7_arsize  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_arvalid (ds7_arvalid ), // (bmc300) => (axi_monitor_s7,axi_slave7,bench)
	.ds7_awaddr  (ds7_awaddr  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awburst (ds7_awburst ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awcache (ds7_awcache ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awid    (ds7_awid    ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awlen   (ds7_awlen   ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awlock  (ds7_awlock  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awprot  (ds7_awprot  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awready (ds7_awready ), // (axi_monitor_s7,bench,bmc300) <= (axi_slave7)
	.ds7_awsize  (ds7_awsize  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_awvalid (ds7_awvalid ), // (bmc300) => (axi_monitor_s7,axi_slave7,bench)
	.ds7_bid     (ds7_bid     ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_bready  (ds7_bready  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_bresp   (ds7_bresp   ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_bvalid  (ds7_bvalid  ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_rdata   (ds7_rdata   ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_rid     (ds7_rid     ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_rlast   (ds7_rlast   ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_rready  (ds7_rready  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_rresp   (ds7_rresp   ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_rvalid  (ds7_rvalid  ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_wdata   (ds7_wdata   ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_wlast   (ds7_wlast   ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_wready  (ds7_wready  ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.ds7_wstrb   (ds7_wstrb   ), // (bmc300) => (axi_monitor_s7,axi_slave7)
	.ds7_wvalid  (ds7_wvalid  ), // (bmc300) => (axi_monitor_s7,axi_slave7)
`endif // ATCBMC300_SLV7_SUPPORT
`ifdef ATCBMC300_SLV8_SUPPORT
	.ds8_araddr  (ds8_araddr  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arburst (ds8_arburst ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arcache (ds8_arcache ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arid    (ds8_arid    ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arlen   (ds8_arlen   ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arlock  (ds8_arlock  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arprot  (ds8_arprot  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arready (ds8_arready ), // (axi_monitor_s8,bench,bmc300) <= (axi_slave8)
	.ds8_arsize  (ds8_arsize  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_arvalid (ds8_arvalid ), // (bmc300) => (axi_monitor_s8,axi_slave8,bench)
	.ds8_awaddr  (ds8_awaddr  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awburst (ds8_awburst ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awcache (ds8_awcache ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awid    (ds8_awid    ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awlen   (ds8_awlen   ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awlock  (ds8_awlock  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awprot  (ds8_awprot  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awready (ds8_awready ), // (axi_monitor_s8,bench,bmc300) <= (axi_slave8)
	.ds8_awsize  (ds8_awsize  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_awvalid (ds8_awvalid ), // (bmc300) => (axi_monitor_s8,axi_slave8,bench)
	.ds8_bid     (ds8_bid     ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_bready  (ds8_bready  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_bresp   (ds8_bresp   ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_bvalid  (ds8_bvalid  ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_rdata   (ds8_rdata   ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_rid     (ds8_rid     ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_rlast   (ds8_rlast   ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_rready  (ds8_rready  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_rresp   (ds8_rresp   ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_rvalid  (ds8_rvalid  ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_wdata   (ds8_wdata   ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_wlast   (ds8_wlast   ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_wready  (ds8_wready  ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.ds8_wstrb   (ds8_wstrb   ), // (bmc300) => (axi_monitor_s8,axi_slave8)
	.ds8_wvalid  (ds8_wvalid  ), // (bmc300) => (axi_monitor_s8,axi_slave8)
`endif // ATCBMC300_SLV8_SUPPORT
`ifdef ATCBMC300_SLV9_SUPPORT
	.ds9_araddr  (ds9_araddr  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arburst (ds9_arburst ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arcache (ds9_arcache ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arid    (ds9_arid    ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arlen   (ds9_arlen   ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arlock  (ds9_arlock  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arprot  (ds9_arprot  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arready (ds9_arready ), // (axi_monitor_s9,bench,bmc300) <= (axi_slave9)
	.ds9_arsize  (ds9_arsize  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_arvalid (ds9_arvalid ), // (bmc300) => (axi_monitor_s9,axi_slave9,bench)
	.ds9_awaddr  (ds9_awaddr  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awburst (ds9_awburst ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awcache (ds9_awcache ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awid    (ds9_awid    ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awlen   (ds9_awlen   ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awlock  (ds9_awlock  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awprot  (ds9_awprot  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awready (ds9_awready ), // (axi_monitor_s9,bench,bmc300) <= (axi_slave9)
	.ds9_awsize  (ds9_awsize  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_awvalid (ds9_awvalid ), // (bmc300) => (axi_monitor_s9,axi_slave9,bench)
	.ds9_bid     (ds9_bid     ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_bready  (ds9_bready  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_bresp   (ds9_bresp   ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_bvalid  (ds9_bvalid  ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_rdata   (ds9_rdata   ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_rid     (ds9_rid     ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_rlast   (ds9_rlast   ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_rready  (ds9_rready  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_rresp   (ds9_rresp   ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_rvalid  (ds9_rvalid  ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_wdata   (ds9_wdata   ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_wlast   (ds9_wlast   ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_wready  (ds9_wready  ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.ds9_wstrb   (ds9_wstrb   ), // (bmc300) => (axi_monitor_s9,axi_slave9)
	.ds9_wvalid  (ds9_wvalid  ), // (bmc300) => (axi_monitor_s9,axi_slave9)
`endif // ATCBMC300_SLV9_SUPPORT
`ifdef ATCBMC300_SLV10_SUPPORT
	.ds10_araddr (ds10_araddr ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arburst(ds10_arburst), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arcache(ds10_arcache), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arid   (ds10_arid   ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arlen  (ds10_arlen  ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arlock (ds10_arlock ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arprot (ds10_arprot ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arready(ds10_arready), // (axi_monitor_s10,bench,bmc300) <= (axi_slave10)
	.ds10_arsize (ds10_arsize ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_arvalid(ds10_arvalid), // (bmc300) => (axi_monitor_s10,axi_slave10,bench)
	.ds10_awaddr (ds10_awaddr ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awburst(ds10_awburst), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awcache(ds10_awcache), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awid   (ds10_awid   ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awlen  (ds10_awlen  ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awlock (ds10_awlock ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awprot (ds10_awprot ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awready(ds10_awready), // (axi_monitor_s10,bench,bmc300) <= (axi_slave10)
	.ds10_awsize (ds10_awsize ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_awvalid(ds10_awvalid), // (bmc300) => (axi_monitor_s10,axi_slave10,bench)
	.ds10_bid    (ds10_bid    ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_bready (ds10_bready ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_bresp  (ds10_bresp  ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_bvalid (ds10_bvalid ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_rdata  (ds10_rdata  ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_rid    (ds10_rid    ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_rlast  (ds10_rlast  ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_rready (ds10_rready ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_rresp  (ds10_rresp  ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_rvalid (ds10_rvalid ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_wdata  (ds10_wdata  ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_wlast  (ds10_wlast  ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_wready (ds10_wready ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.ds10_wstrb  (ds10_wstrb  ), // (bmc300) => (axi_monitor_s10,axi_slave10)
	.ds10_wvalid (ds10_wvalid ), // (bmc300) => (axi_monitor_s10,axi_slave10)
`endif // ATCBMC300_SLV10_SUPPORT
`ifdef ATCBMC300_SLV11_SUPPORT
	.ds11_araddr (ds11_araddr ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arburst(ds11_arburst), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arcache(ds11_arcache), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arid   (ds11_arid   ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arlen  (ds11_arlen  ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arlock (ds11_arlock ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arprot (ds11_arprot ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arready(ds11_arready), // (axi_monitor_s11,bench,bmc300) <= (axi_slave11)
	.ds11_arsize (ds11_arsize ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_arvalid(ds11_arvalid), // (bmc300) => (axi_monitor_s11,axi_slave11,bench)
	.ds11_awaddr (ds11_awaddr ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awburst(ds11_awburst), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awcache(ds11_awcache), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awid   (ds11_awid   ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awlen  (ds11_awlen  ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awlock (ds11_awlock ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awprot (ds11_awprot ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awready(ds11_awready), // (axi_monitor_s11,bench,bmc300) <= (axi_slave11)
	.ds11_awsize (ds11_awsize ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_awvalid(ds11_awvalid), // (bmc300) => (axi_monitor_s11,axi_slave11,bench)
	.ds11_bid    (ds11_bid    ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_bready (ds11_bready ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_bresp  (ds11_bresp  ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_bvalid (ds11_bvalid ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_rdata  (ds11_rdata  ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_rid    (ds11_rid    ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_rlast  (ds11_rlast  ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_rready (ds11_rready ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_rresp  (ds11_rresp  ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_rvalid (ds11_rvalid ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_wdata  (ds11_wdata  ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_wlast  (ds11_wlast  ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_wready (ds11_wready ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.ds11_wstrb  (ds11_wstrb  ), // (bmc300) => (axi_monitor_s11,axi_slave11)
	.ds11_wvalid (ds11_wvalid ), // (bmc300) => (axi_monitor_s11,axi_slave11)
`endif // ATCBMC300_SLV11_SUPPORT
`ifdef ATCBMC300_SLV12_SUPPORT
	.ds12_araddr (ds12_araddr ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arburst(ds12_arburst), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arcache(ds12_arcache), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arid   (ds12_arid   ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arlen  (ds12_arlen  ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arlock (ds12_arlock ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arprot (ds12_arprot ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arready(ds12_arready), // (axi_monitor_s12,bench,bmc300) <= (axi_slave12)
	.ds12_arsize (ds12_arsize ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_arvalid(ds12_arvalid), // (bmc300) => (axi_monitor_s12,axi_slave12,bench)
	.ds12_awaddr (ds12_awaddr ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awburst(ds12_awburst), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awcache(ds12_awcache), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awid   (ds12_awid   ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awlen  (ds12_awlen  ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awlock (ds12_awlock ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awprot (ds12_awprot ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awready(ds12_awready), // (axi_monitor_s12,bench,bmc300) <= (axi_slave12)
	.ds12_awsize (ds12_awsize ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_awvalid(ds12_awvalid), // (bmc300) => (axi_monitor_s12,axi_slave12,bench)
	.ds12_bid    (ds12_bid    ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_bready (ds12_bready ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_bresp  (ds12_bresp  ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_bvalid (ds12_bvalid ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_rdata  (ds12_rdata  ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_rid    (ds12_rid    ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_rlast  (ds12_rlast  ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_rready (ds12_rready ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_rresp  (ds12_rresp  ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_rvalid (ds12_rvalid ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_wdata  (ds12_wdata  ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_wlast  (ds12_wlast  ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_wready (ds12_wready ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.ds12_wstrb  (ds12_wstrb  ), // (bmc300) => (axi_monitor_s12,axi_slave12)
	.ds12_wvalid (ds12_wvalid ), // (bmc300) => (axi_monitor_s12,axi_slave12)
`endif // ATCBMC300_SLV12_SUPPORT
`ifdef ATCBMC300_SLV13_SUPPORT
	.ds13_araddr (ds13_araddr ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arburst(ds13_arburst), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arcache(ds13_arcache), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arid   (ds13_arid   ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arlen  (ds13_arlen  ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arlock (ds13_arlock ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arprot (ds13_arprot ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arready(ds13_arready), // (axi_monitor_s13,bench,bmc300) <= (axi_slave13)
	.ds13_arsize (ds13_arsize ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_arvalid(ds13_arvalid), // (bmc300) => (axi_monitor_s13,axi_slave13,bench)
	.ds13_awaddr (ds13_awaddr ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awburst(ds13_awburst), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awcache(ds13_awcache), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awid   (ds13_awid   ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awlen  (ds13_awlen  ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awlock (ds13_awlock ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awprot (ds13_awprot ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awready(ds13_awready), // (axi_monitor_s13,bench,bmc300) <= (axi_slave13)
	.ds13_awsize (ds13_awsize ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_awvalid(ds13_awvalid), // (bmc300) => (axi_monitor_s13,axi_slave13,bench)
	.ds13_bid    (ds13_bid    ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_bready (ds13_bready ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_bresp  (ds13_bresp  ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_bvalid (ds13_bvalid ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_rdata  (ds13_rdata  ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_rid    (ds13_rid    ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_rlast  (ds13_rlast  ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_rready (ds13_rready ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_rresp  (ds13_rresp  ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_rvalid (ds13_rvalid ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_wdata  (ds13_wdata  ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_wlast  (ds13_wlast  ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_wready (ds13_wready ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.ds13_wstrb  (ds13_wstrb  ), // (bmc300) => (axi_monitor_s13,axi_slave13)
	.ds13_wvalid (ds13_wvalid ), // (bmc300) => (axi_monitor_s13,axi_slave13)
`endif // ATCBMC300_SLV13_SUPPORT
`ifdef ATCBMC300_SLV14_SUPPORT
	.ds14_araddr (ds14_araddr ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arburst(ds14_arburst), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arcache(ds14_arcache), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arid   (ds14_arid   ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arlen  (ds14_arlen  ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arlock (ds14_arlock ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arprot (ds14_arprot ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arready(ds14_arready), // (axi_monitor_s14,bench,bmc300) <= (axi_slave14)
	.ds14_arsize (ds14_arsize ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_arvalid(ds14_arvalid), // (bmc300) => (axi_monitor_s14,axi_slave14,bench)
	.ds14_awaddr (ds14_awaddr ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awburst(ds14_awburst), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awcache(ds14_awcache), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awid   (ds14_awid   ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awlen  (ds14_awlen  ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awlock (ds14_awlock ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awprot (ds14_awprot ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awready(ds14_awready), // (axi_monitor_s14,bench,bmc300) <= (axi_slave14)
	.ds14_awsize (ds14_awsize ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_awvalid(ds14_awvalid), // (bmc300) => (axi_monitor_s14,axi_slave14,bench)
	.ds14_bid    (ds14_bid    ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_bready (ds14_bready ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_bresp  (ds14_bresp  ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_bvalid (ds14_bvalid ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_rdata  (ds14_rdata  ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_rid    (ds14_rid    ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_rlast  (ds14_rlast  ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_rready (ds14_rready ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_rresp  (ds14_rresp  ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_rvalid (ds14_rvalid ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_wdata  (ds14_wdata  ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_wlast  (ds14_wlast  ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_wready (ds14_wready ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.ds14_wstrb  (ds14_wstrb  ), // (bmc300) => (axi_monitor_s14,axi_slave14)
	.ds14_wvalid (ds14_wvalid ), // (bmc300) => (axi_monitor_s14,axi_slave14)
`endif // ATCBMC300_SLV14_SUPPORT
`ifdef ATCBMC300_SLV15_SUPPORT
	.ds15_araddr (ds15_araddr ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arburst(ds15_arburst), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arcache(ds15_arcache), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arid   (ds15_arid   ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arlen  (ds15_arlen  ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arlock (ds15_arlock ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arprot (ds15_arprot ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arready(ds15_arready), // (axi_monitor_s15,bench,bmc300) <= (axi_slave15)
	.ds15_arsize (ds15_arsize ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_arvalid(ds15_arvalid), // (bmc300) => (axi_monitor_s15,axi_slave15,bench)
	.ds15_awaddr (ds15_awaddr ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awburst(ds15_awburst), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awcache(ds15_awcache), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awid   (ds15_awid   ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awlen  (ds15_awlen  ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awlock (ds15_awlock ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awprot (ds15_awprot ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awready(ds15_awready), // (axi_monitor_s15,bench,bmc300) <= (axi_slave15)
	.ds15_awsize (ds15_awsize ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_awvalid(ds15_awvalid), // (bmc300) => (axi_monitor_s15,axi_slave15,bench)
	.ds15_bid    (ds15_bid    ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_bready (ds15_bready ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_bresp  (ds15_bresp  ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_bvalid (ds15_bvalid ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_rdata  (ds15_rdata  ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_rid    (ds15_rid    ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_rlast  (ds15_rlast  ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_rready (ds15_rready ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_rresp  (ds15_rresp  ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_rvalid (ds15_rvalid ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_wdata  (ds15_wdata  ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_wlast  (ds15_wlast  ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_wready (ds15_wready ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.ds15_wstrb  (ds15_wstrb  ), // (bmc300) => (axi_monitor_s15,axi_slave15)
	.ds15_wvalid (ds15_wvalid ), // (bmc300) => (axi_monitor_s15,axi_slave15)
`endif // ATCBMC300_SLV15_SUPPORT
`ifdef ATCBMC300_SLV16_SUPPORT
	.ds16_araddr (ds16_araddr ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arburst(ds16_arburst), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arcache(ds16_arcache), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arid   (ds16_arid   ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arlen  (ds16_arlen  ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arlock (ds16_arlock ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arprot (ds16_arprot ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arready(ds16_arready), // (axi_monitor_s16,bench,bmc300) <= (axi_slave16)
	.ds16_arsize (ds16_arsize ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_arvalid(ds16_arvalid), // (bmc300) => (axi_monitor_s16,axi_slave16,bench)
	.ds16_awaddr (ds16_awaddr ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awburst(ds16_awburst), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awcache(ds16_awcache), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awid   (ds16_awid   ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awlen  (ds16_awlen  ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awlock (ds16_awlock ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awprot (ds16_awprot ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awready(ds16_awready), // (axi_monitor_s16,bench,bmc300) <= (axi_slave16)
	.ds16_awsize (ds16_awsize ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_awvalid(ds16_awvalid), // (bmc300) => (axi_monitor_s16,axi_slave16,bench)
	.ds16_bid    (ds16_bid    ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_bready (ds16_bready ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_bresp  (ds16_bresp  ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_bvalid (ds16_bvalid ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_rdata  (ds16_rdata  ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_rid    (ds16_rid    ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_rlast  (ds16_rlast  ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_rready (ds16_rready ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_rresp  (ds16_rresp  ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_rvalid (ds16_rvalid ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_wdata  (ds16_wdata  ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_wlast  (ds16_wlast  ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_wready (ds16_wready ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.ds16_wstrb  (ds16_wstrb  ), // (bmc300) => (axi_monitor_s16,axi_slave16)
	.ds16_wvalid (ds16_wvalid ), // (bmc300) => (axi_monitor_s16,axi_slave16)
`endif // ATCBMC300_SLV16_SUPPORT
`ifdef ATCBMC300_SLV17_SUPPORT
	.ds17_araddr (ds17_araddr ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arburst(ds17_arburst), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arcache(ds17_arcache), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arid   (ds17_arid   ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arlen  (ds17_arlen  ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arlock (ds17_arlock ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arprot (ds17_arprot ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arready(ds17_arready), // (axi_monitor_s17,bench,bmc300) <= (axi_slave17)
	.ds17_arsize (ds17_arsize ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_arvalid(ds17_arvalid), // (bmc300) => (axi_monitor_s17,axi_slave17,bench)
	.ds17_awaddr (ds17_awaddr ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awburst(ds17_awburst), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awcache(ds17_awcache), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awid   (ds17_awid   ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awlen  (ds17_awlen  ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awlock (ds17_awlock ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awprot (ds17_awprot ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awready(ds17_awready), // (axi_monitor_s17,bench,bmc300) <= (axi_slave17)
	.ds17_awsize (ds17_awsize ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_awvalid(ds17_awvalid), // (bmc300) => (axi_monitor_s17,axi_slave17,bench)
	.ds17_bid    (ds17_bid    ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_bready (ds17_bready ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_bresp  (ds17_bresp  ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_bvalid (ds17_bvalid ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_rdata  (ds17_rdata  ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_rid    (ds17_rid    ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_rlast  (ds17_rlast  ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_rready (ds17_rready ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_rresp  (ds17_rresp  ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_rvalid (ds17_rvalid ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_wdata  (ds17_wdata  ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_wlast  (ds17_wlast  ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_wready (ds17_wready ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.ds17_wstrb  (ds17_wstrb  ), // (bmc300) => (axi_monitor_s17,axi_slave17)
	.ds17_wvalid (ds17_wvalid ), // (bmc300) => (axi_monitor_s17,axi_slave17)
`endif // ATCBMC300_SLV17_SUPPORT
`ifdef ATCBMC300_SLV18_SUPPORT
	.ds18_araddr (ds18_araddr ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arburst(ds18_arburst), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arcache(ds18_arcache), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arid   (ds18_arid   ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arlen  (ds18_arlen  ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arlock (ds18_arlock ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arprot (ds18_arprot ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arready(ds18_arready), // (axi_monitor_s18,bench,bmc300) <= (axi_slave18)
	.ds18_arsize (ds18_arsize ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_arvalid(ds18_arvalid), // (bmc300) => (axi_monitor_s18,axi_slave18,bench)
	.ds18_awaddr (ds18_awaddr ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awburst(ds18_awburst), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awcache(ds18_awcache), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awid   (ds18_awid   ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awlen  (ds18_awlen  ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awlock (ds18_awlock ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awprot (ds18_awprot ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awready(ds18_awready), // (axi_monitor_s18,bench,bmc300) <= (axi_slave18)
	.ds18_awsize (ds18_awsize ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_awvalid(ds18_awvalid), // (bmc300) => (axi_monitor_s18,axi_slave18,bench)
	.ds18_bid    (ds18_bid    ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_bready (ds18_bready ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_bresp  (ds18_bresp  ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_bvalid (ds18_bvalid ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_rdata  (ds18_rdata  ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_rid    (ds18_rid    ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_rlast  (ds18_rlast  ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_rready (ds18_rready ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_rresp  (ds18_rresp  ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_rvalid (ds18_rvalid ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_wdata  (ds18_wdata  ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_wlast  (ds18_wlast  ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_wready (ds18_wready ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.ds18_wstrb  (ds18_wstrb  ), // (bmc300) => (axi_monitor_s18,axi_slave18)
	.ds18_wvalid (ds18_wvalid ), // (bmc300) => (axi_monitor_s18,axi_slave18)
`endif // ATCBMC300_SLV18_SUPPORT
`ifdef ATCBMC300_SLV19_SUPPORT
	.ds19_araddr (ds19_araddr ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arburst(ds19_arburst), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arcache(ds19_arcache), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arid   (ds19_arid   ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arlen  (ds19_arlen  ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arlock (ds19_arlock ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arprot (ds19_arprot ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arready(ds19_arready), // (axi_monitor_s19,bench,bmc300) <= (axi_slave19)
	.ds19_arsize (ds19_arsize ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_arvalid(ds19_arvalid), // (bmc300) => (axi_monitor_s19,axi_slave19,bench)
	.ds19_awaddr (ds19_awaddr ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awburst(ds19_awburst), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awcache(ds19_awcache), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awid   (ds19_awid   ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awlen  (ds19_awlen  ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awlock (ds19_awlock ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awprot (ds19_awprot ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awready(ds19_awready), // (axi_monitor_s19,bench,bmc300) <= (axi_slave19)
	.ds19_awsize (ds19_awsize ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_awvalid(ds19_awvalid), // (bmc300) => (axi_monitor_s19,axi_slave19,bench)
	.ds19_bid    (ds19_bid    ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_bready (ds19_bready ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_bresp  (ds19_bresp  ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_bvalid (ds19_bvalid ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_rdata  (ds19_rdata  ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_rid    (ds19_rid    ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_rlast  (ds19_rlast  ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_rready (ds19_rready ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_rresp  (ds19_rresp  ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_rvalid (ds19_rvalid ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_wdata  (ds19_wdata  ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_wlast  (ds19_wlast  ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_wready (ds19_wready ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.ds19_wstrb  (ds19_wstrb  ), // (bmc300) => (axi_monitor_s19,axi_slave19)
	.ds19_wvalid (ds19_wvalid ), // (bmc300) => (axi_monitor_s19,axi_slave19)
`endif // ATCBMC300_SLV19_SUPPORT
`ifdef ATCBMC300_SLV20_SUPPORT
	.ds20_araddr (ds20_araddr ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arburst(ds20_arburst), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arcache(ds20_arcache), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arid   (ds20_arid   ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arlen  (ds20_arlen  ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arlock (ds20_arlock ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arprot (ds20_arprot ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arready(ds20_arready), // (axi_monitor_s20,bench,bmc300) <= (axi_slave20)
	.ds20_arsize (ds20_arsize ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_arvalid(ds20_arvalid), // (bmc300) => (axi_monitor_s20,axi_slave20,bench)
	.ds20_awaddr (ds20_awaddr ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awburst(ds20_awburst), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awcache(ds20_awcache), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awid   (ds20_awid   ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awlen  (ds20_awlen  ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awlock (ds20_awlock ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awprot (ds20_awprot ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awready(ds20_awready), // (axi_monitor_s20,bench,bmc300) <= (axi_slave20)
	.ds20_awsize (ds20_awsize ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_awvalid(ds20_awvalid), // (bmc300) => (axi_monitor_s20,axi_slave20,bench)
	.ds20_bid    (ds20_bid    ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_bready (ds20_bready ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_bresp  (ds20_bresp  ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_bvalid (ds20_bvalid ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_rdata  (ds20_rdata  ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_rid    (ds20_rid    ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_rlast  (ds20_rlast  ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_rready (ds20_rready ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_rresp  (ds20_rresp  ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_rvalid (ds20_rvalid ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_wdata  (ds20_wdata  ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_wlast  (ds20_wlast  ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_wready (ds20_wready ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.ds20_wstrb  (ds20_wstrb  ), // (bmc300) => (axi_monitor_s20,axi_slave20)
	.ds20_wvalid (ds20_wvalid ), // (bmc300) => (axi_monitor_s20,axi_slave20)
`endif // ATCBMC300_SLV20_SUPPORT
`ifdef ATCBMC300_SLV21_SUPPORT
	.ds21_araddr (ds21_araddr ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arburst(ds21_arburst), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arcache(ds21_arcache), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arid   (ds21_arid   ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arlen  (ds21_arlen  ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arlock (ds21_arlock ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arprot (ds21_arprot ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arready(ds21_arready), // (axi_monitor_s21,bench,bmc300) <= (axi_slave21)
	.ds21_arsize (ds21_arsize ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_arvalid(ds21_arvalid), // (bmc300) => (axi_monitor_s21,axi_slave21,bench)
	.ds21_awaddr (ds21_awaddr ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awburst(ds21_awburst), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awcache(ds21_awcache), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awid   (ds21_awid   ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awlen  (ds21_awlen  ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awlock (ds21_awlock ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awprot (ds21_awprot ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awready(ds21_awready), // (axi_monitor_s21,bench,bmc300) <= (axi_slave21)
	.ds21_awsize (ds21_awsize ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_awvalid(ds21_awvalid), // (bmc300) => (axi_monitor_s21,axi_slave21,bench)
	.ds21_bid    (ds21_bid    ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_bready (ds21_bready ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_bresp  (ds21_bresp  ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_bvalid (ds21_bvalid ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_rdata  (ds21_rdata  ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_rid    (ds21_rid    ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_rlast  (ds21_rlast  ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_rready (ds21_rready ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_rresp  (ds21_rresp  ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_rvalid (ds21_rvalid ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_wdata  (ds21_wdata  ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_wlast  (ds21_wlast  ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_wready (ds21_wready ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.ds21_wstrb  (ds21_wstrb  ), // (bmc300) => (axi_monitor_s21,axi_slave21)
	.ds21_wvalid (ds21_wvalid ), // (bmc300) => (axi_monitor_s21,axi_slave21)
`endif // ATCBMC300_SLV21_SUPPORT
`ifdef ATCBMC300_SLV22_SUPPORT
	.ds22_araddr (ds22_araddr ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arburst(ds22_arburst), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arcache(ds22_arcache), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arid   (ds22_arid   ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arlen  (ds22_arlen  ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arlock (ds22_arlock ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arprot (ds22_arprot ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arready(ds22_arready), // (axi_monitor_s22,bench,bmc300) <= (axi_slave22)
	.ds22_arsize (ds22_arsize ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_arvalid(ds22_arvalid), // (bmc300) => (axi_monitor_s22,axi_slave22,bench)
	.ds22_awaddr (ds22_awaddr ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awburst(ds22_awburst), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awcache(ds22_awcache), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awid   (ds22_awid   ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awlen  (ds22_awlen  ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awlock (ds22_awlock ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awprot (ds22_awprot ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awready(ds22_awready), // (axi_monitor_s22,bench,bmc300) <= (axi_slave22)
	.ds22_awsize (ds22_awsize ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_awvalid(ds22_awvalid), // (bmc300) => (axi_monitor_s22,axi_slave22,bench)
	.ds22_bid    (ds22_bid    ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_bready (ds22_bready ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_bresp  (ds22_bresp  ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_bvalid (ds22_bvalid ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_rdata  (ds22_rdata  ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_rid    (ds22_rid    ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_rlast  (ds22_rlast  ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_rready (ds22_rready ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_rresp  (ds22_rresp  ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_rvalid (ds22_rvalid ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_wdata  (ds22_wdata  ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_wlast  (ds22_wlast  ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_wready (ds22_wready ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.ds22_wstrb  (ds22_wstrb  ), // (bmc300) => (axi_monitor_s22,axi_slave22)
	.ds22_wvalid (ds22_wvalid ), // (bmc300) => (axi_monitor_s22,axi_slave22)
`endif // ATCBMC300_SLV22_SUPPORT
`ifdef ATCBMC300_SLV23_SUPPORT
	.ds23_araddr (ds23_araddr ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arburst(ds23_arburst), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arcache(ds23_arcache), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arid   (ds23_arid   ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arlen  (ds23_arlen  ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arlock (ds23_arlock ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arprot (ds23_arprot ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arready(ds23_arready), // (axi_monitor_s23,bench,bmc300) <= (axi_slave23)
	.ds23_arsize (ds23_arsize ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_arvalid(ds23_arvalid), // (bmc300) => (axi_monitor_s23,axi_slave23,bench)
	.ds23_awaddr (ds23_awaddr ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awburst(ds23_awburst), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awcache(ds23_awcache), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awid   (ds23_awid   ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awlen  (ds23_awlen  ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awlock (ds23_awlock ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awprot (ds23_awprot ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awready(ds23_awready), // (axi_monitor_s23,bench,bmc300) <= (axi_slave23)
	.ds23_awsize (ds23_awsize ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_awvalid(ds23_awvalid), // (bmc300) => (axi_monitor_s23,axi_slave23,bench)
	.ds23_bid    (ds23_bid    ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_bready (ds23_bready ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_bresp  (ds23_bresp  ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_bvalid (ds23_bvalid ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_rdata  (ds23_rdata  ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_rid    (ds23_rid    ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_rlast  (ds23_rlast  ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_rready (ds23_rready ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_rresp  (ds23_rresp  ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_rvalid (ds23_rvalid ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_wdata  (ds23_wdata  ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_wlast  (ds23_wlast  ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_wready (ds23_wready ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.ds23_wstrb  (ds23_wstrb  ), // (bmc300) => (axi_monitor_s23,axi_slave23)
	.ds23_wvalid (ds23_wvalid ), // (bmc300) => (axi_monitor_s23,axi_slave23)
`endif // ATCBMC300_SLV23_SUPPORT
`ifdef ATCBMC300_SLV24_SUPPORT
	.ds24_araddr (ds24_araddr ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arburst(ds24_arburst), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arcache(ds24_arcache), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arid   (ds24_arid   ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arlen  (ds24_arlen  ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arlock (ds24_arlock ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arprot (ds24_arprot ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arready(ds24_arready), // (axi_monitor_s24,bench,bmc300) <= (axi_slave24)
	.ds24_arsize (ds24_arsize ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_arvalid(ds24_arvalid), // (bmc300) => (axi_monitor_s24,axi_slave24,bench)
	.ds24_awaddr (ds24_awaddr ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awburst(ds24_awburst), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awcache(ds24_awcache), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awid   (ds24_awid   ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awlen  (ds24_awlen  ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awlock (ds24_awlock ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awprot (ds24_awprot ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awready(ds24_awready), // (axi_monitor_s24,bench,bmc300) <= (axi_slave24)
	.ds24_awsize (ds24_awsize ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_awvalid(ds24_awvalid), // (bmc300) => (axi_monitor_s24,axi_slave24,bench)
	.ds24_bid    (ds24_bid    ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_bready (ds24_bready ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_bresp  (ds24_bresp  ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_bvalid (ds24_bvalid ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_rdata  (ds24_rdata  ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_rid    (ds24_rid    ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_rlast  (ds24_rlast  ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_rready (ds24_rready ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_rresp  (ds24_rresp  ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_rvalid (ds24_rvalid ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_wdata  (ds24_wdata  ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_wlast  (ds24_wlast  ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_wready (ds24_wready ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.ds24_wstrb  (ds24_wstrb  ), // (bmc300) => (axi_monitor_s24,axi_slave24)
	.ds24_wvalid (ds24_wvalid ), // (bmc300) => (axi_monitor_s24,axi_slave24)
`endif // ATCBMC300_SLV24_SUPPORT
`ifdef ATCBMC300_SLV25_SUPPORT
	.ds25_araddr (ds25_araddr ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arburst(ds25_arburst), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arcache(ds25_arcache), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arid   (ds25_arid   ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arlen  (ds25_arlen  ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arlock (ds25_arlock ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arprot (ds25_arprot ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arready(ds25_arready), // (axi_monitor_s25,bench,bmc300) <= (axi_slave25)
	.ds25_arsize (ds25_arsize ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_arvalid(ds25_arvalid), // (bmc300) => (axi_monitor_s25,axi_slave25,bench)
	.ds25_awaddr (ds25_awaddr ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awburst(ds25_awburst), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awcache(ds25_awcache), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awid   (ds25_awid   ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awlen  (ds25_awlen  ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awlock (ds25_awlock ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awprot (ds25_awprot ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awready(ds25_awready), // (axi_monitor_s25,bench,bmc300) <= (axi_slave25)
	.ds25_awsize (ds25_awsize ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_awvalid(ds25_awvalid), // (bmc300) => (axi_monitor_s25,axi_slave25,bench)
	.ds25_bid    (ds25_bid    ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_bready (ds25_bready ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_bresp  (ds25_bresp  ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_bvalid (ds25_bvalid ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_rdata  (ds25_rdata  ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_rid    (ds25_rid    ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_rlast  (ds25_rlast  ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_rready (ds25_rready ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_rresp  (ds25_rresp  ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_rvalid (ds25_rvalid ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_wdata  (ds25_wdata  ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_wlast  (ds25_wlast  ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_wready (ds25_wready ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.ds25_wstrb  (ds25_wstrb  ), // (bmc300) => (axi_monitor_s25,axi_slave25)
	.ds25_wvalid (ds25_wvalid ), // (bmc300) => (axi_monitor_s25,axi_slave25)
`endif // ATCBMC300_SLV25_SUPPORT
`ifdef ATCBMC300_SLV26_SUPPORT
	.ds26_araddr (ds26_araddr ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arburst(ds26_arburst), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arcache(ds26_arcache), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arid   (ds26_arid   ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arlen  (ds26_arlen  ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arlock (ds26_arlock ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arprot (ds26_arprot ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arready(ds26_arready), // (axi_monitor_s26,bench,bmc300) <= (axi_slave26)
	.ds26_arsize (ds26_arsize ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_arvalid(ds26_arvalid), // (bmc300) => (axi_monitor_s26,axi_slave26,bench)
	.ds26_awaddr (ds26_awaddr ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awburst(ds26_awburst), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awcache(ds26_awcache), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awid   (ds26_awid   ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awlen  (ds26_awlen  ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awlock (ds26_awlock ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awprot (ds26_awprot ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awready(ds26_awready), // (axi_monitor_s26,bench,bmc300) <= (axi_slave26)
	.ds26_awsize (ds26_awsize ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_awvalid(ds26_awvalid), // (bmc300) => (axi_monitor_s26,axi_slave26,bench)
	.ds26_bid    (ds26_bid    ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_bready (ds26_bready ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_bresp  (ds26_bresp  ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_bvalid (ds26_bvalid ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_rdata  (ds26_rdata  ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_rid    (ds26_rid    ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_rlast  (ds26_rlast  ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_rready (ds26_rready ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_rresp  (ds26_rresp  ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_rvalid (ds26_rvalid ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_wdata  (ds26_wdata  ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_wlast  (ds26_wlast  ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_wready (ds26_wready ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.ds26_wstrb  (ds26_wstrb  ), // (bmc300) => (axi_monitor_s26,axi_slave26)
	.ds26_wvalid (ds26_wvalid ), // (bmc300) => (axi_monitor_s26,axi_slave26)
`endif // ATCBMC300_SLV26_SUPPORT
`ifdef ATCBMC300_SLV27_SUPPORT
	.ds27_araddr (ds27_araddr ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arburst(ds27_arburst), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arcache(ds27_arcache), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arid   (ds27_arid   ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arlen  (ds27_arlen  ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arlock (ds27_arlock ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arprot (ds27_arprot ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arready(ds27_arready), // (axi_monitor_s27,bench,bmc300) <= (axi_slave27)
	.ds27_arsize (ds27_arsize ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_arvalid(ds27_arvalid), // (bmc300) => (axi_monitor_s27,axi_slave27,bench)
	.ds27_awaddr (ds27_awaddr ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awburst(ds27_awburst), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awcache(ds27_awcache), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awid   (ds27_awid   ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awlen  (ds27_awlen  ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awlock (ds27_awlock ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awprot (ds27_awprot ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awready(ds27_awready), // (axi_monitor_s27,bench,bmc300) <= (axi_slave27)
	.ds27_awsize (ds27_awsize ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_awvalid(ds27_awvalid), // (bmc300) => (axi_monitor_s27,axi_slave27,bench)
	.ds27_bid    (ds27_bid    ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_bready (ds27_bready ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_bresp  (ds27_bresp  ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_bvalid (ds27_bvalid ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_rdata  (ds27_rdata  ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_rid    (ds27_rid    ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_rlast  (ds27_rlast  ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_rready (ds27_rready ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_rresp  (ds27_rresp  ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_rvalid (ds27_rvalid ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_wdata  (ds27_wdata  ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_wlast  (ds27_wlast  ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_wready (ds27_wready ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.ds27_wstrb  (ds27_wstrb  ), // (bmc300) => (axi_monitor_s27,axi_slave27)
	.ds27_wvalid (ds27_wvalid ), // (bmc300) => (axi_monitor_s27,axi_slave27)
`endif // ATCBMC300_SLV27_SUPPORT
`ifdef ATCBMC300_SLV28_SUPPORT
	.ds28_araddr (ds28_araddr ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arburst(ds28_arburst), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arcache(ds28_arcache), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arid   (ds28_arid   ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arlen  (ds28_arlen  ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arlock (ds28_arlock ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arprot (ds28_arprot ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arready(ds28_arready), // (axi_monitor_s28,bench,bmc300) <= (axi_slave28)
	.ds28_arsize (ds28_arsize ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_arvalid(ds28_arvalid), // (bmc300) => (axi_monitor_s28,axi_slave28,bench)
	.ds28_awaddr (ds28_awaddr ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awburst(ds28_awburst), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awcache(ds28_awcache), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awid   (ds28_awid   ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awlen  (ds28_awlen  ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awlock (ds28_awlock ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awprot (ds28_awprot ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awready(ds28_awready), // (axi_monitor_s28,bench,bmc300) <= (axi_slave28)
	.ds28_awsize (ds28_awsize ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_awvalid(ds28_awvalid), // (bmc300) => (axi_monitor_s28,axi_slave28,bench)
	.ds28_bid    (ds28_bid    ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_bready (ds28_bready ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_bresp  (ds28_bresp  ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_bvalid (ds28_bvalid ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_rdata  (ds28_rdata  ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_rid    (ds28_rid    ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_rlast  (ds28_rlast  ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_rready (ds28_rready ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_rresp  (ds28_rresp  ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_rvalid (ds28_rvalid ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_wdata  (ds28_wdata  ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_wlast  (ds28_wlast  ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_wready (ds28_wready ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.ds28_wstrb  (ds28_wstrb  ), // (bmc300) => (axi_monitor_s28,axi_slave28)
	.ds28_wvalid (ds28_wvalid ), // (bmc300) => (axi_monitor_s28,axi_slave28)
`endif // ATCBMC300_SLV28_SUPPORT
`ifdef ATCBMC300_SLV29_SUPPORT
	.ds29_araddr (ds29_araddr ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arburst(ds29_arburst), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arcache(ds29_arcache), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arid   (ds29_arid   ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arlen  (ds29_arlen  ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arlock (ds29_arlock ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arprot (ds29_arprot ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arready(ds29_arready), // (axi_monitor_s29,bench,bmc300) <= (axi_slave29)
	.ds29_arsize (ds29_arsize ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_arvalid(ds29_arvalid), // (bmc300) => (axi_monitor_s29,axi_slave29,bench)
	.ds29_awaddr (ds29_awaddr ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awburst(ds29_awburst), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awcache(ds29_awcache), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awid   (ds29_awid   ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awlen  (ds29_awlen  ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awlock (ds29_awlock ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awprot (ds29_awprot ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awready(ds29_awready), // (axi_monitor_s29,bench,bmc300) <= (axi_slave29)
	.ds29_awsize (ds29_awsize ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_awvalid(ds29_awvalid), // (bmc300) => (axi_monitor_s29,axi_slave29,bench)
	.ds29_bid    (ds29_bid    ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_bready (ds29_bready ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_bresp  (ds29_bresp  ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_bvalid (ds29_bvalid ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_rdata  (ds29_rdata  ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_rid    (ds29_rid    ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_rlast  (ds29_rlast  ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_rready (ds29_rready ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_rresp  (ds29_rresp  ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_rvalid (ds29_rvalid ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_wdata  (ds29_wdata  ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_wlast  (ds29_wlast  ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_wready (ds29_wready ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.ds29_wstrb  (ds29_wstrb  ), // (bmc300) => (axi_monitor_s29,axi_slave29)
	.ds29_wvalid (ds29_wvalid ), // (bmc300) => (axi_monitor_s29,axi_slave29)
`endif // ATCBMC300_SLV29_SUPPORT
`ifdef ATCBMC300_SLV30_SUPPORT
	.ds30_araddr (ds30_araddr ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arburst(ds30_arburst), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arcache(ds30_arcache), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arid   (ds30_arid   ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arlen  (ds30_arlen  ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arlock (ds30_arlock ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arprot (ds30_arprot ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arready(ds30_arready), // (axi_monitor_s30,bench,bmc300) <= (axi_slave30)
	.ds30_arsize (ds30_arsize ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_arvalid(ds30_arvalid), // (bmc300) => (axi_monitor_s30,axi_slave30,bench)
	.ds30_awaddr (ds30_awaddr ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awburst(ds30_awburst), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awcache(ds30_awcache), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awid   (ds30_awid   ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awlen  (ds30_awlen  ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awlock (ds30_awlock ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awprot (ds30_awprot ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awready(ds30_awready), // (axi_monitor_s30,bench,bmc300) <= (axi_slave30)
	.ds30_awsize (ds30_awsize ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_awvalid(ds30_awvalid), // (bmc300) => (axi_monitor_s30,axi_slave30,bench)
	.ds30_bid    (ds30_bid    ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_bready (ds30_bready ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_bresp  (ds30_bresp  ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_bvalid (ds30_bvalid ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_rdata  (ds30_rdata  ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_rid    (ds30_rid    ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_rlast  (ds30_rlast  ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_rready (ds30_rready ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_rresp  (ds30_rresp  ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_rvalid (ds30_rvalid ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_wdata  (ds30_wdata  ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_wlast  (ds30_wlast  ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_wready (ds30_wready ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.ds30_wstrb  (ds30_wstrb  ), // (bmc300) => (axi_monitor_s30,axi_slave30)
	.ds30_wvalid (ds30_wvalid ), // (bmc300) => (axi_monitor_s30,axi_slave30)
`endif // ATCBMC300_SLV30_SUPPORT
`ifdef ATCBMC300_SLV31_SUPPORT
	.ds31_araddr (ds31_araddr ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arburst(ds31_arburst), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arcache(ds31_arcache), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arid   (ds31_arid   ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arlen  (ds31_arlen  ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arlock (ds31_arlock ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arprot (ds31_arprot ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arready(ds31_arready), // (axi_monitor_s31,bench,bmc300) <= (axi_slave31)
	.ds31_arsize (ds31_arsize ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_arvalid(ds31_arvalid), // (bmc300) => (axi_monitor_s31,axi_slave31,bench)
	.ds31_awaddr (ds31_awaddr ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awburst(ds31_awburst), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awcache(ds31_awcache), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awid   (ds31_awid   ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awlen  (ds31_awlen  ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awlock (ds31_awlock ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awprot (ds31_awprot ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awready(ds31_awready), // (axi_monitor_s31,bench,bmc300) <= (axi_slave31)
	.ds31_awsize (ds31_awsize ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_awvalid(ds31_awvalid), // (bmc300) => (axi_monitor_s31,axi_slave31,bench)
	.ds31_bid    (ds31_bid    ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_bready (ds31_bready ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_bresp  (ds31_bresp  ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_bvalid (ds31_bvalid ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_rdata  (ds31_rdata  ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_rid    (ds31_rid    ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_rlast  (ds31_rlast  ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_rready (ds31_rready ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_rresp  (ds31_rresp  ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_rvalid (ds31_rvalid ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_wdata  (ds31_wdata  ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_wlast  (ds31_wlast  ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_wready (ds31_wready ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.ds31_wstrb  (ds31_wstrb  ), // (bmc300) => (axi_monitor_s31,axi_slave31)
	.ds31_wvalid (ds31_wvalid ), // (bmc300) => (axi_monitor_s31,axi_slave31)
`endif // ATCBMC300_SLV31_SUPPORT
`ifdef ATCBMC300_MST1_SUPPORT
	.us1_araddr  (us1_araddr  ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_arburst (us1_arburst ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arcache (us1_arcache ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arid    (us1_arid    ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arlen   (us1_arlen   ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arlock  (us1_arlock  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arprot  (us1_arprot  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arready (us1_arready ), // (bmc300) => (axi_master1,axi_monitor_m1,bench)
	.us1_arsize  (us1_arsize  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_arvalid (us1_arvalid ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_awaddr  (us1_awaddr  ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_awburst (us1_awburst ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awcache (us1_awcache ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awid    (us1_awid    ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awlen   (us1_awlen   ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awlock  (us1_awlock  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awprot  (us1_awprot  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awready (us1_awready ), // (bmc300) => (axi_master1,axi_monitor_m1,bench)
	.us1_awsize  (us1_awsize  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_awvalid (us1_awvalid ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_bid     (us1_bid     ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_bready  (us1_bready  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_bresp   (us1_bresp   ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_bvalid  (us1_bvalid  ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_rdata   (us1_rdata   ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_rid     (us1_rid     ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_rlast   (us1_rlast   ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_rready  (us1_rready  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_rresp   (us1_rresp   ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_rvalid  (us1_rvalid  ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_wdata   (us1_wdata   ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_wlast   (us1_wlast   ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_wready  (us1_wready  ), // (bmc300) => (axi_master1,axi_monitor_m1)
	.us1_wstrb   (us1_wstrb   ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.us1_wvalid  (us1_wvalid  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
`endif // ATCBMC300_MST1_SUPPORT
`ifdef ATCBMC300_MST2_SUPPORT
	.us2_araddr  (us2_araddr  ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_arburst (us2_arburst ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arcache (us2_arcache ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arid    (us2_arid    ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arlen   (us2_arlen   ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arlock  (us2_arlock  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arprot  (us2_arprot  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arready (us2_arready ), // (bmc300) => (axi_master2,axi_monitor_m2,bench)
	.us2_arsize  (us2_arsize  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_arvalid (us2_arvalid ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_awaddr  (us2_awaddr  ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_awburst (us2_awburst ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awcache (us2_awcache ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awid    (us2_awid    ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awlen   (us2_awlen   ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awlock  (us2_awlock  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awprot  (us2_awprot  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awready (us2_awready ), // (bmc300) => (axi_master2,axi_monitor_m2,bench)
	.us2_awsize  (us2_awsize  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_awvalid (us2_awvalid ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_bid     (us2_bid     ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_bready  (us2_bready  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_bresp   (us2_bresp   ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_bvalid  (us2_bvalid  ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_rdata   (us2_rdata   ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_rid     (us2_rid     ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_rlast   (us2_rlast   ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_rready  (us2_rready  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_rresp   (us2_rresp   ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_rvalid  (us2_rvalid  ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_wdata   (us2_wdata   ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_wlast   (us2_wlast   ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_wready  (us2_wready  ), // (bmc300) => (axi_master2,axi_monitor_m2)
	.us2_wstrb   (us2_wstrb   ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.us2_wvalid  (us2_wvalid  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
`endif // ATCBMC300_MST2_SUPPORT
`ifdef ATCBMC300_MST3_SUPPORT
	.us3_araddr  (us3_araddr  ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_arburst (us3_arburst ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arcache (us3_arcache ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arid    (us3_arid    ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arlen   (us3_arlen   ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arlock  (us3_arlock  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arprot  (us3_arprot  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arready (us3_arready ), // (bmc300) => (axi_master3,axi_monitor_m3,bench)
	.us3_arsize  (us3_arsize  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_arvalid (us3_arvalid ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_awaddr  (us3_awaddr  ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_awburst (us3_awburst ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awcache (us3_awcache ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awid    (us3_awid    ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awlen   (us3_awlen   ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awlock  (us3_awlock  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awprot  (us3_awprot  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awready (us3_awready ), // (bmc300) => (axi_master3,axi_monitor_m3,bench)
	.us3_awsize  (us3_awsize  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_awvalid (us3_awvalid ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_bid     (us3_bid     ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_bready  (us3_bready  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_bresp   (us3_bresp   ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_bvalid  (us3_bvalid  ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_rdata   (us3_rdata   ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_rid     (us3_rid     ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_rlast   (us3_rlast   ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_rready  (us3_rready  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_rresp   (us3_rresp   ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_rvalid  (us3_rvalid  ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_wdata   (us3_wdata   ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_wlast   (us3_wlast   ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_wready  (us3_wready  ), // (bmc300) => (axi_master3,axi_monitor_m3)
	.us3_wstrb   (us3_wstrb   ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.us3_wvalid  (us3_wvalid  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
`endif // ATCBMC300_MST3_SUPPORT
`ifdef ATCBMC300_MST4_SUPPORT
	.us4_araddr  (us4_araddr  ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_arburst (us4_arburst ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arcache (us4_arcache ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arid    (us4_arid    ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arlen   (us4_arlen   ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arlock  (us4_arlock  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arprot  (us4_arprot  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arready (us4_arready ), // (bmc300) => (axi_master4,axi_monitor_m4,bench)
	.us4_arsize  (us4_arsize  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_arvalid (us4_arvalid ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_awaddr  (us4_awaddr  ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_awburst (us4_awburst ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awcache (us4_awcache ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awid    (us4_awid    ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awlen   (us4_awlen   ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awlock  (us4_awlock  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awprot  (us4_awprot  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awready (us4_awready ), // (bmc300) => (axi_master4,axi_monitor_m4,bench)
	.us4_awsize  (us4_awsize  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_awvalid (us4_awvalid ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_bid     (us4_bid     ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_bready  (us4_bready  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_bresp   (us4_bresp   ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_bvalid  (us4_bvalid  ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_rdata   (us4_rdata   ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_rid     (us4_rid     ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_rlast   (us4_rlast   ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_rready  (us4_rready  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_rresp   (us4_rresp   ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_rvalid  (us4_rvalid  ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_wdata   (us4_wdata   ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_wlast   (us4_wlast   ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_wready  (us4_wready  ), // (bmc300) => (axi_master4,axi_monitor_m4)
	.us4_wstrb   (us4_wstrb   ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.us4_wvalid  (us4_wvalid  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
`endif // ATCBMC300_MST4_SUPPORT
`ifdef ATCBMC300_MST5_SUPPORT
	.us5_araddr  (us5_araddr  ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_arburst (us5_arburst ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arcache (us5_arcache ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arid    (us5_arid    ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arlen   (us5_arlen   ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arlock  (us5_arlock  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arprot  (us5_arprot  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arready (us5_arready ), // (bmc300) => (axi_master5,axi_monitor_m5,bench)
	.us5_arsize  (us5_arsize  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_arvalid (us5_arvalid ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_awaddr  (us5_awaddr  ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_awburst (us5_awburst ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awcache (us5_awcache ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awid    (us5_awid    ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awlen   (us5_awlen   ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awlock  (us5_awlock  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awprot  (us5_awprot  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awready (us5_awready ), // (bmc300) => (axi_master5,axi_monitor_m5,bench)
	.us5_awsize  (us5_awsize  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_awvalid (us5_awvalid ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_bid     (us5_bid     ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_bready  (us5_bready  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_bresp   (us5_bresp   ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_bvalid  (us5_bvalid  ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_rdata   (us5_rdata   ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_rid     (us5_rid     ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_rlast   (us5_rlast   ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_rready  (us5_rready  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_rresp   (us5_rresp   ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_rvalid  (us5_rvalid  ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_wdata   (us5_wdata   ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_wlast   (us5_wlast   ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_wready  (us5_wready  ), // (bmc300) => (axi_master5,axi_monitor_m5)
	.us5_wstrb   (us5_wstrb   ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.us5_wvalid  (us5_wvalid  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
`endif // ATCBMC300_MST5_SUPPORT
`ifdef ATCBMC300_MST6_SUPPORT
	.us6_araddr  (us6_araddr  ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_arburst (us6_arburst ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arcache (us6_arcache ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arid    (us6_arid    ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arlen   (us6_arlen   ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arlock  (us6_arlock  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arprot  (us6_arprot  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arready (us6_arready ), // (bmc300) => (axi_master6,axi_monitor_m6,bench)
	.us6_arsize  (us6_arsize  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_arvalid (us6_arvalid ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_awaddr  (us6_awaddr  ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_awburst (us6_awburst ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awcache (us6_awcache ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awid    (us6_awid    ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awlen   (us6_awlen   ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awlock  (us6_awlock  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awprot  (us6_awprot  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awready (us6_awready ), // (bmc300) => (axi_master6,axi_monitor_m6,bench)
	.us6_awsize  (us6_awsize  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_awvalid (us6_awvalid ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_bid     (us6_bid     ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_bready  (us6_bready  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_bresp   (us6_bresp   ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_bvalid  (us6_bvalid  ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_rdata   (us6_rdata   ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_rid     (us6_rid     ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_rlast   (us6_rlast   ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_rready  (us6_rready  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_rresp   (us6_rresp   ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_rvalid  (us6_rvalid  ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_wdata   (us6_wdata   ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_wlast   (us6_wlast   ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_wready  (us6_wready  ), // (bmc300) => (axi_master6,axi_monitor_m6)
	.us6_wstrb   (us6_wstrb   ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.us6_wvalid  (us6_wvalid  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
`endif // ATCBMC300_MST6_SUPPORT
`ifdef ATCBMC300_MST7_SUPPORT
	.us7_araddr  (us7_araddr  ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_arburst (us7_arburst ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arcache (us7_arcache ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arid    (us7_arid    ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arlen   (us7_arlen   ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arlock  (us7_arlock  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arprot  (us7_arprot  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arready (us7_arready ), // (bmc300) => (axi_master7,axi_monitor_m7,bench)
	.us7_arsize  (us7_arsize  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_arvalid (us7_arvalid ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_awaddr  (us7_awaddr  ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_awburst (us7_awburst ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awcache (us7_awcache ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awid    (us7_awid    ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awlen   (us7_awlen   ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awlock  (us7_awlock  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awprot  (us7_awprot  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awready (us7_awready ), // (bmc300) => (axi_master7,axi_monitor_m7,bench)
	.us7_awsize  (us7_awsize  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_awvalid (us7_awvalid ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_bid     (us7_bid     ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_bready  (us7_bready  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_bresp   (us7_bresp   ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_bvalid  (us7_bvalid  ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_rdata   (us7_rdata   ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_rid     (us7_rid     ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_rlast   (us7_rlast   ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_rready  (us7_rready  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_rresp   (us7_rresp   ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_rvalid  (us7_rvalid  ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_wdata   (us7_wdata   ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_wlast   (us7_wlast   ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_wready  (us7_wready  ), // (bmc300) => (axi_master7,axi_monitor_m7)
	.us7_wstrb   (us7_wstrb   ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.us7_wvalid  (us7_wvalid  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
`endif // ATCBMC300_MST7_SUPPORT
`ifdef ATCBMC300_MST8_SUPPORT
	.us8_araddr  (us8_araddr  ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_arburst (us8_arburst ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arcache (us8_arcache ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arid    (us8_arid    ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arlen   (us8_arlen   ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arlock  (us8_arlock  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arprot  (us8_arprot  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arready (us8_arready ), // (bmc300) => (axi_master8,axi_monitor_m8,bench)
	.us8_arsize  (us8_arsize  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_arvalid (us8_arvalid ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_awaddr  (us8_awaddr  ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_awburst (us8_awburst ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awcache (us8_awcache ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awid    (us8_awid    ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awlen   (us8_awlen   ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awlock  (us8_awlock  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awprot  (us8_awprot  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awready (us8_awready ), // (bmc300) => (axi_master8,axi_monitor_m8,bench)
	.us8_awsize  (us8_awsize  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_awvalid (us8_awvalid ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_bid     (us8_bid     ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_bready  (us8_bready  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_bresp   (us8_bresp   ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_bvalid  (us8_bvalid  ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_rdata   (us8_rdata   ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_rid     (us8_rid     ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_rlast   (us8_rlast   ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_rready  (us8_rready  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_rresp   (us8_rresp   ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_rvalid  (us8_rvalid  ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_wdata   (us8_wdata   ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_wlast   (us8_wlast   ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_wready  (us8_wready  ), // (bmc300) => (axi_master8,axi_monitor_m8)
	.us8_wstrb   (us8_wstrb   ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.us8_wvalid  (us8_wvalid  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
`endif // ATCBMC300_MST8_SUPPORT
`ifdef ATCBMC300_MST9_SUPPORT
	.us9_araddr  (us9_araddr  ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_arburst (us9_arburst ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arcache (us9_arcache ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arid    (us9_arid    ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arlen   (us9_arlen   ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arlock  (us9_arlock  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arprot  (us9_arprot  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arready (us9_arready ), // (bmc300) => (axi_master9,axi_monitor_m9,bench)
	.us9_arsize  (us9_arsize  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_arvalid (us9_arvalid ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_awaddr  (us9_awaddr  ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_awburst (us9_awburst ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awcache (us9_awcache ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awid    (us9_awid    ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awlen   (us9_awlen   ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awlock  (us9_awlock  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awprot  (us9_awprot  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awready (us9_awready ), // (bmc300) => (axi_master9,axi_monitor_m9,bench)
	.us9_awsize  (us9_awsize  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_awvalid (us9_awvalid ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_bid     (us9_bid     ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_bready  (us9_bready  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_bresp   (us9_bresp   ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_bvalid  (us9_bvalid  ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_rdata   (us9_rdata   ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_rid     (us9_rid     ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_rlast   (us9_rlast   ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_rready  (us9_rready  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_rresp   (us9_rresp   ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_rvalid  (us9_rvalid  ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_wdata   (us9_wdata   ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_wlast   (us9_wlast   ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_wready  (us9_wready  ), // (bmc300) => (axi_master9,axi_monitor_m9)
	.us9_wstrb   (us9_wstrb   ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.us9_wvalid  (us9_wvalid  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
`endif // ATCBMC300_MST9_SUPPORT
`ifdef ATCBMC300_MST10_SUPPORT
	.us10_araddr (us10_araddr ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_arburst(us10_arburst), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arcache(us10_arcache), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arid   (us10_arid   ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arlen  (us10_arlen  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arlock (us10_arlock ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arprot (us10_arprot ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arready(us10_arready), // (bmc300) => (axi_master10,axi_monitor_m10,bench)
	.us10_arsize (us10_arsize ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_arvalid(us10_arvalid), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_awaddr (us10_awaddr ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_awburst(us10_awburst), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awcache(us10_awcache), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awid   (us10_awid   ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awlen  (us10_awlen  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awlock (us10_awlock ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awprot (us10_awprot ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awready(us10_awready), // (bmc300) => (axi_master10,axi_monitor_m10,bench)
	.us10_awsize (us10_awsize ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_awvalid(us10_awvalid), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_bid    (us10_bid    ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_bready (us10_bready ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_bresp  (us10_bresp  ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_bvalid (us10_bvalid ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_rdata  (us10_rdata  ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_rid    (us10_rid    ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_rlast  (us10_rlast  ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_rready (us10_rready ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_rresp  (us10_rresp  ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_rvalid (us10_rvalid ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_wdata  (us10_wdata  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_wlast  (us10_wlast  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_wready (us10_wready ), // (bmc300) => (axi_master10,axi_monitor_m10)
	.us10_wstrb  (us10_wstrb  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.us10_wvalid (us10_wvalid ), // (axi_monitor_m10,bmc300) <= (axi_master10)
`endif // ATCBMC300_MST10_SUPPORT
`ifdef ATCBMC300_MST11_SUPPORT
	.us11_araddr (us11_araddr ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_arburst(us11_arburst), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arcache(us11_arcache), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arid   (us11_arid   ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arlen  (us11_arlen  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arlock (us11_arlock ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arprot (us11_arprot ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arready(us11_arready), // (bmc300) => (axi_master11,axi_monitor_m11,bench)
	.us11_arsize (us11_arsize ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_arvalid(us11_arvalid), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_awaddr (us11_awaddr ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_awburst(us11_awburst), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awcache(us11_awcache), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awid   (us11_awid   ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awlen  (us11_awlen  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awlock (us11_awlock ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awprot (us11_awprot ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awready(us11_awready), // (bmc300) => (axi_master11,axi_monitor_m11,bench)
	.us11_awsize (us11_awsize ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_awvalid(us11_awvalid), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_bid    (us11_bid    ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_bready (us11_bready ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_bresp  (us11_bresp  ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_bvalid (us11_bvalid ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_rdata  (us11_rdata  ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_rid    (us11_rid    ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_rlast  (us11_rlast  ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_rready (us11_rready ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_rresp  (us11_rresp  ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_rvalid (us11_rvalid ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_wdata  (us11_wdata  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_wlast  (us11_wlast  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_wready (us11_wready ), // (bmc300) => (axi_master11,axi_monitor_m11)
	.us11_wstrb  (us11_wstrb  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.us11_wvalid (us11_wvalid ), // (axi_monitor_m11,bmc300) <= (axi_master11)
`endif // ATCBMC300_MST11_SUPPORT
`ifdef ATCBMC300_MST12_SUPPORT
	.us12_araddr (us12_araddr ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_arburst(us12_arburst), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arcache(us12_arcache), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arid   (us12_arid   ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arlen  (us12_arlen  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arlock (us12_arlock ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arprot (us12_arprot ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arready(us12_arready), // (bmc300) => (axi_master12,axi_monitor_m12,bench)
	.us12_arsize (us12_arsize ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_arvalid(us12_arvalid), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_awaddr (us12_awaddr ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_awburst(us12_awburst), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awcache(us12_awcache), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awid   (us12_awid   ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awlen  (us12_awlen  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awlock (us12_awlock ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awprot (us12_awprot ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awready(us12_awready), // (bmc300) => (axi_master12,axi_monitor_m12,bench)
	.us12_awsize (us12_awsize ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_awvalid(us12_awvalid), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_bid    (us12_bid    ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_bready (us12_bready ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_bresp  (us12_bresp  ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_bvalid (us12_bvalid ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_rdata  (us12_rdata  ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_rid    (us12_rid    ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_rlast  (us12_rlast  ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_rready (us12_rready ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_rresp  (us12_rresp  ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_rvalid (us12_rvalid ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_wdata  (us12_wdata  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_wlast  (us12_wlast  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_wready (us12_wready ), // (bmc300) => (axi_master12,axi_monitor_m12)
	.us12_wstrb  (us12_wstrb  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.us12_wvalid (us12_wvalid ), // (axi_monitor_m12,bmc300) <= (axi_master12)
`endif // ATCBMC300_MST12_SUPPORT
`ifdef ATCBMC300_MST13_SUPPORT
	.us13_araddr (us13_araddr ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_arburst(us13_arburst), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arcache(us13_arcache), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arid   (us13_arid   ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arlen  (us13_arlen  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arlock (us13_arlock ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arprot (us13_arprot ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arready(us13_arready), // (bmc300) => (axi_master13,axi_monitor_m13,bench)
	.us13_arsize (us13_arsize ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_arvalid(us13_arvalid), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_awaddr (us13_awaddr ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_awburst(us13_awburst), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awcache(us13_awcache), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awid   (us13_awid   ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awlen  (us13_awlen  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awlock (us13_awlock ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awprot (us13_awprot ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awready(us13_awready), // (bmc300) => (axi_master13,axi_monitor_m13,bench)
	.us13_awsize (us13_awsize ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_awvalid(us13_awvalid), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_bid    (us13_bid    ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_bready (us13_bready ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_bresp  (us13_bresp  ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_bvalid (us13_bvalid ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_rdata  (us13_rdata  ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_rid    (us13_rid    ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_rlast  (us13_rlast  ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_rready (us13_rready ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_rresp  (us13_rresp  ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_rvalid (us13_rvalid ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_wdata  (us13_wdata  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_wlast  (us13_wlast  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_wready (us13_wready ), // (bmc300) => (axi_master13,axi_monitor_m13)
	.us13_wstrb  (us13_wstrb  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.us13_wvalid (us13_wvalid ), // (axi_monitor_m13,bmc300) <= (axi_master13)
`endif // ATCBMC300_MST13_SUPPORT
`ifdef ATCBMC300_MST14_SUPPORT
	.us14_araddr (us14_araddr ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_arburst(us14_arburst), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arcache(us14_arcache), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arid   (us14_arid   ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arlen  (us14_arlen  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arlock (us14_arlock ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arprot (us14_arprot ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arready(us14_arready), // (bmc300) => (axi_master14,axi_monitor_m14,bench)
	.us14_arsize (us14_arsize ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_arvalid(us14_arvalid), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_awaddr (us14_awaddr ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_awburst(us14_awburst), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awcache(us14_awcache), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awid   (us14_awid   ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awlen  (us14_awlen  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awlock (us14_awlock ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awprot (us14_awprot ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awready(us14_awready), // (bmc300) => (axi_master14,axi_monitor_m14,bench)
	.us14_awsize (us14_awsize ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_awvalid(us14_awvalid), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_bid    (us14_bid    ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_bready (us14_bready ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_bresp  (us14_bresp  ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_bvalid (us14_bvalid ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_rdata  (us14_rdata  ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_rid    (us14_rid    ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_rlast  (us14_rlast  ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_rready (us14_rready ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_rresp  (us14_rresp  ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_rvalid (us14_rvalid ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_wdata  (us14_wdata  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_wlast  (us14_wlast  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_wready (us14_wready ), // (bmc300) => (axi_master14,axi_monitor_m14)
	.us14_wstrb  (us14_wstrb  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.us14_wvalid (us14_wvalid ), // (axi_monitor_m14,bmc300) <= (axi_master14)
`endif // ATCBMC300_MST14_SUPPORT
`ifdef ATCBMC300_MST15_SUPPORT
	.us15_araddr (us15_araddr ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_arburst(us15_arburst), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arcache(us15_arcache), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arid   (us15_arid   ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arlen  (us15_arlen  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arlock (us15_arlock ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arprot (us15_arprot ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arready(us15_arready), // (bmc300) => (axi_master15,axi_monitor_m15,bench)
	.us15_arsize (us15_arsize ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_arvalid(us15_arvalid), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_awaddr (us15_awaddr ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_awburst(us15_awburst), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awcache(us15_awcache), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awid   (us15_awid   ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awlen  (us15_awlen  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awlock (us15_awlock ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awprot (us15_awprot ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awready(us15_awready), // (bmc300) => (axi_master15,axi_monitor_m15,bench)
	.us15_awsize (us15_awsize ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_awvalid(us15_awvalid), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_bid    (us15_bid    ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_bready (us15_bready ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_bresp  (us15_bresp  ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_bvalid (us15_bvalid ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_rdata  (us15_rdata  ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_rid    (us15_rid    ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_rlast  (us15_rlast  ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_rready (us15_rready ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_rresp  (us15_rresp  ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_rvalid (us15_rvalid ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_wdata  (us15_wdata  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_wlast  (us15_wlast  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_wready (us15_wready ), // (bmc300) => (axi_master15,axi_monitor_m15)
	.us15_wstrb  (us15_wstrb  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.us15_wvalid (us15_wvalid ), // (axi_monitor_m15,bmc300) <= (axi_master15)
`endif // ATCBMC300_MST15_SUPPORT
	.aclk        (aclk        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn     (aresetn     )  // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
); // end of bmc300

defparam bench.ADDR_WIDTH = ADDR_WIDTH;
defparam bench.DATA_SIZE = DATA_SIZE;
defparam bench.DS_ID_WIDTH = DS_ID_WIDTH;
defparam bench.ERROR_PROBABILITY = `NDS_ERROR_PROBABILITY;
blk_tb bench (
`ifdef ATCBMC300_MST0_SUPPORT
	.us0_arvalid (us0_arvalid ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_arready (us0_arready ), // (axi_master0,axi_monitor_m0,bench) <= (bmc300)
	.us0_araddr  (us0_araddr  ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_awvalid (us0_awvalid ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.us0_awready (us0_awready ), // (axi_master0,axi_monitor_m0,bench) <= (bmc300)
	.us0_awaddr  (us0_awaddr  ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
`endif // ATCBMC300_MST0_SUPPORT
`ifdef ATCBMC300_MST1_SUPPORT
	.us1_arvalid (us1_arvalid ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_arready (us1_arready ), // (axi_master1,axi_monitor_m1,bench) <= (bmc300)
	.us1_araddr  (us1_araddr  ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_awvalid (us1_awvalid ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.us1_awready (us1_awready ), // (axi_master1,axi_monitor_m1,bench) <= (bmc300)
	.us1_awaddr  (us1_awaddr  ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
`endif // ATCBMC300_MST1_SUPPORT
`ifdef ATCBMC300_MST2_SUPPORT
	.us2_arvalid (us2_arvalid ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_arready (us2_arready ), // (axi_master2,axi_monitor_m2,bench) <= (bmc300)
	.us2_araddr  (us2_araddr  ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_awvalid (us2_awvalid ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.us2_awready (us2_awready ), // (axi_master2,axi_monitor_m2,bench) <= (bmc300)
	.us2_awaddr  (us2_awaddr  ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
`endif // ATCBMC300_MST2_SUPPORT
`ifdef ATCBMC300_MST3_SUPPORT
	.us3_arvalid (us3_arvalid ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_arready (us3_arready ), // (axi_master3,axi_monitor_m3,bench) <= (bmc300)
	.us3_araddr  (us3_araddr  ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_awvalid (us3_awvalid ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.us3_awready (us3_awready ), // (axi_master3,axi_monitor_m3,bench) <= (bmc300)
	.us3_awaddr  (us3_awaddr  ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
`endif // ATCBMC300_MST3_SUPPORT
`ifdef ATCBMC300_MST4_SUPPORT
	.us4_arvalid (us4_arvalid ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_arready (us4_arready ), // (axi_master4,axi_monitor_m4,bench) <= (bmc300)
	.us4_araddr  (us4_araddr  ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_awvalid (us4_awvalid ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.us4_awready (us4_awready ), // (axi_master4,axi_monitor_m4,bench) <= (bmc300)
	.us4_awaddr  (us4_awaddr  ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
`endif // ATCBMC300_MST4_SUPPORT
`ifdef ATCBMC300_MST5_SUPPORT
	.us5_arvalid (us5_arvalid ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_arready (us5_arready ), // (axi_master5,axi_monitor_m5,bench) <= (bmc300)
	.us5_araddr  (us5_araddr  ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_awvalid (us5_awvalid ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.us5_awready (us5_awready ), // (axi_master5,axi_monitor_m5,bench) <= (bmc300)
	.us5_awaddr  (us5_awaddr  ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
`endif // ATCBMC300_MST5_SUPPORT
`ifdef ATCBMC300_MST6_SUPPORT
	.us6_arvalid (us6_arvalid ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_arready (us6_arready ), // (axi_master6,axi_monitor_m6,bench) <= (bmc300)
	.us6_araddr  (us6_araddr  ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_awvalid (us6_awvalid ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.us6_awready (us6_awready ), // (axi_master6,axi_monitor_m6,bench) <= (bmc300)
	.us6_awaddr  (us6_awaddr  ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
`endif // ATCBMC300_MST6_SUPPORT
`ifdef ATCBMC300_MST7_SUPPORT
	.us7_arvalid (us7_arvalid ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_arready (us7_arready ), // (axi_master7,axi_monitor_m7,bench) <= (bmc300)
	.us7_araddr  (us7_araddr  ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_awvalid (us7_awvalid ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.us7_awready (us7_awready ), // (axi_master7,axi_monitor_m7,bench) <= (bmc300)
	.us7_awaddr  (us7_awaddr  ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
`endif // ATCBMC300_MST7_SUPPORT
`ifdef ATCBMC300_MST8_SUPPORT
	.us8_arvalid (us8_arvalid ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_arready (us8_arready ), // (axi_master8,axi_monitor_m8,bench) <= (bmc300)
	.us8_araddr  (us8_araddr  ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_awvalid (us8_awvalid ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.us8_awready (us8_awready ), // (axi_master8,axi_monitor_m8,bench) <= (bmc300)
	.us8_awaddr  (us8_awaddr  ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
`endif // ATCBMC300_MST8_SUPPORT
`ifdef ATCBMC300_MST9_SUPPORT
	.us9_arvalid (us9_arvalid ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_arready (us9_arready ), // (axi_master9,axi_monitor_m9,bench) <= (bmc300)
	.us9_araddr  (us9_araddr  ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_awvalid (us9_awvalid ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.us9_awready (us9_awready ), // (axi_master9,axi_monitor_m9,bench) <= (bmc300)
	.us9_awaddr  (us9_awaddr  ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
`endif // ATCBMC300_MST9_SUPPORT
`ifdef ATCBMC300_MST10_SUPPORT
	.us10_arvalid(us10_arvalid), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_arready(us10_arready), // (axi_master10,axi_monitor_m10,bench) <= (bmc300)
	.us10_araddr (us10_araddr ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_awvalid(us10_awvalid), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.us10_awready(us10_awready), // (axi_master10,axi_monitor_m10,bench) <= (bmc300)
	.us10_awaddr (us10_awaddr ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
`endif // ATCBMC300_MST10_SUPPORT
`ifdef ATCBMC300_MST11_SUPPORT
	.us11_arvalid(us11_arvalid), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_arready(us11_arready), // (axi_master11,axi_monitor_m11,bench) <= (bmc300)
	.us11_araddr (us11_araddr ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_awvalid(us11_awvalid), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.us11_awready(us11_awready), // (axi_master11,axi_monitor_m11,bench) <= (bmc300)
	.us11_awaddr (us11_awaddr ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
`endif // ATCBMC300_MST11_SUPPORT
`ifdef ATCBMC300_MST12_SUPPORT
	.us12_arvalid(us12_arvalid), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_arready(us12_arready), // (axi_master12,axi_monitor_m12,bench) <= (bmc300)
	.us12_araddr (us12_araddr ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_awvalid(us12_awvalid), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.us12_awready(us12_awready), // (axi_master12,axi_monitor_m12,bench) <= (bmc300)
	.us12_awaddr (us12_awaddr ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
`endif // ATCBMC300_MST12_SUPPORT
`ifdef ATCBMC300_MST13_SUPPORT
	.us13_arvalid(us13_arvalid), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_arready(us13_arready), // (axi_master13,axi_monitor_m13,bench) <= (bmc300)
	.us13_araddr (us13_araddr ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_awvalid(us13_awvalid), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.us13_awready(us13_awready), // (axi_master13,axi_monitor_m13,bench) <= (bmc300)
	.us13_awaddr (us13_awaddr ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
`endif // ATCBMC300_MST13_SUPPORT
`ifdef ATCBMC300_MST14_SUPPORT
	.us14_arvalid(us14_arvalid), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_arready(us14_arready), // (axi_master14,axi_monitor_m14,bench) <= (bmc300)
	.us14_araddr (us14_araddr ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_awvalid(us14_awvalid), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.us14_awready(us14_awready), // (axi_master14,axi_monitor_m14,bench) <= (bmc300)
	.us14_awaddr (us14_awaddr ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
`endif // ATCBMC300_MST14_SUPPORT
`ifdef ATCBMC300_MST15_SUPPORT
	.us15_arvalid(us15_arvalid), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_arready(us15_arready), // (axi_master15,axi_monitor_m15,bench) <= (bmc300)
	.us15_araddr (us15_araddr ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_awvalid(us15_awvalid), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.us15_awready(us15_awready), // (axi_master15,axi_monitor_m15,bench) <= (bmc300)
	.us15_awaddr (us15_awaddr ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
`endif // ATCBMC300_MST15_SUPPORT
`ifdef ATCBMC300_SLV1_SUPPORT
	.ds1_arvalid (ds1_arvalid ), // (axi_monitor_s1,axi_slave1,bench) <= (bmc300)
	.ds1_arready (ds1_arready ), // (axi_monitor_s1,bench,bmc300) <= (axi_slave1)
	.ds1_awvalid (ds1_awvalid ), // (axi_monitor_s1,axi_slave1,bench) <= (bmc300)
	.ds1_awready (ds1_awready ), // (axi_monitor_s1,bench,bmc300) <= (axi_slave1)
`endif // ATCBMC300_SLV1_SUPPORT
`ifdef ATCBMC300_SLV2_SUPPORT
	.ds2_arvalid (ds2_arvalid ), // (axi_monitor_s2,axi_slave2,bench) <= (bmc300)
	.ds2_arready (ds2_arready ), // (axi_monitor_s2,bench,bmc300) <= (axi_slave2)
	.ds2_awvalid (ds2_awvalid ), // (axi_monitor_s2,axi_slave2,bench) <= (bmc300)
	.ds2_awready (ds2_awready ), // (axi_monitor_s2,bench,bmc300) <= (axi_slave2)
`endif // ATCBMC300_SLV2_SUPPORT
`ifdef ATCBMC300_SLV3_SUPPORT
	.ds3_arvalid (ds3_arvalid ), // (axi_monitor_s3,axi_slave3,bench) <= (bmc300)
	.ds3_arready (ds3_arready ), // (axi_monitor_s3,bench,bmc300) <= (axi_slave3)
	.ds3_awvalid (ds3_awvalid ), // (axi_monitor_s3,axi_slave3,bench) <= (bmc300)
	.ds3_awready (ds3_awready ), // (axi_monitor_s3,bench,bmc300) <= (axi_slave3)
`endif // ATCBMC300_SLV3_SUPPORT
`ifdef ATCBMC300_SLV4_SUPPORT
	.ds4_arvalid (ds4_arvalid ), // (axi_monitor_s4,axi_slave4,bench) <= (bmc300)
	.ds4_arready (ds4_arready ), // (axi_monitor_s4,bench,bmc300) <= (axi_slave4)
	.ds4_awvalid (ds4_awvalid ), // (axi_monitor_s4,axi_slave4,bench) <= (bmc300)
	.ds4_awready (ds4_awready ), // (axi_monitor_s4,bench,bmc300) <= (axi_slave4)
`endif // ATCBMC300_SLV4_SUPPORT
`ifdef ATCBMC300_SLV5_SUPPORT
	.ds5_arvalid (ds5_arvalid ), // (axi_monitor_s5,axi_slave5,bench) <= (bmc300)
	.ds5_arready (ds5_arready ), // (axi_monitor_s5,bench,bmc300) <= (axi_slave5)
	.ds5_awvalid (ds5_awvalid ), // (axi_monitor_s5,axi_slave5,bench) <= (bmc300)
	.ds5_awready (ds5_awready ), // (axi_monitor_s5,bench,bmc300) <= (axi_slave5)
`endif // ATCBMC300_SLV5_SUPPORT
`ifdef ATCBMC300_SLV6_SUPPORT
	.ds6_arvalid (ds6_arvalid ), // (axi_monitor_s6,axi_slave6,bench) <= (bmc300)
	.ds6_arready (ds6_arready ), // (axi_monitor_s6,bench,bmc300) <= (axi_slave6)
	.ds6_awvalid (ds6_awvalid ), // (axi_monitor_s6,axi_slave6,bench) <= (bmc300)
	.ds6_awready (ds6_awready ), // (axi_monitor_s6,bench,bmc300) <= (axi_slave6)
`endif // ATCBMC300_SLV6_SUPPORT
`ifdef ATCBMC300_SLV7_SUPPORT
	.ds7_arvalid (ds7_arvalid ), // (axi_monitor_s7,axi_slave7,bench) <= (bmc300)
	.ds7_arready (ds7_arready ), // (axi_monitor_s7,bench,bmc300) <= (axi_slave7)
	.ds7_awvalid (ds7_awvalid ), // (axi_monitor_s7,axi_slave7,bench) <= (bmc300)
	.ds7_awready (ds7_awready ), // (axi_monitor_s7,bench,bmc300) <= (axi_slave7)
`endif // ATCBMC300_SLV7_SUPPORT
`ifdef ATCBMC300_SLV8_SUPPORT
	.ds8_arvalid (ds8_arvalid ), // (axi_monitor_s8,axi_slave8,bench) <= (bmc300)
	.ds8_arready (ds8_arready ), // (axi_monitor_s8,bench,bmc300) <= (axi_slave8)
	.ds8_awvalid (ds8_awvalid ), // (axi_monitor_s8,axi_slave8,bench) <= (bmc300)
	.ds8_awready (ds8_awready ), // (axi_monitor_s8,bench,bmc300) <= (axi_slave8)
`endif // ATCBMC300_SLV8_SUPPORT
`ifdef ATCBMC300_SLV9_SUPPORT
	.ds9_arvalid (ds9_arvalid ), // (axi_monitor_s9,axi_slave9,bench) <= (bmc300)
	.ds9_arready (ds9_arready ), // (axi_monitor_s9,bench,bmc300) <= (axi_slave9)
	.ds9_awvalid (ds9_awvalid ), // (axi_monitor_s9,axi_slave9,bench) <= (bmc300)
	.ds9_awready (ds9_awready ), // (axi_monitor_s9,bench,bmc300) <= (axi_slave9)
`endif // ATCBMC300_SLV9_SUPPORT
`ifdef ATCBMC300_SLV10_SUPPORT
	.ds10_arvalid(ds10_arvalid), // (axi_monitor_s10,axi_slave10,bench) <= (bmc300)
	.ds10_arready(ds10_arready), // (axi_monitor_s10,bench,bmc300) <= (axi_slave10)
	.ds10_awvalid(ds10_awvalid), // (axi_monitor_s10,axi_slave10,bench) <= (bmc300)
	.ds10_awready(ds10_awready), // (axi_monitor_s10,bench,bmc300) <= (axi_slave10)
`endif // ATCBMC300_SLV10_SUPPORT
`ifdef ATCBMC300_SLV11_SUPPORT
	.ds11_arvalid(ds11_arvalid), // (axi_monitor_s11,axi_slave11,bench) <= (bmc300)
	.ds11_arready(ds11_arready), // (axi_monitor_s11,bench,bmc300) <= (axi_slave11)
	.ds11_awvalid(ds11_awvalid), // (axi_monitor_s11,axi_slave11,bench) <= (bmc300)
	.ds11_awready(ds11_awready), // (axi_monitor_s11,bench,bmc300) <= (axi_slave11)
`endif // ATCBMC300_SLV11_SUPPORT
`ifdef ATCBMC300_SLV12_SUPPORT
	.ds12_arvalid(ds12_arvalid), // (axi_monitor_s12,axi_slave12,bench) <= (bmc300)
	.ds12_arready(ds12_arready), // (axi_monitor_s12,bench,bmc300) <= (axi_slave12)
	.ds12_awvalid(ds12_awvalid), // (axi_monitor_s12,axi_slave12,bench) <= (bmc300)
	.ds12_awready(ds12_awready), // (axi_monitor_s12,bench,bmc300) <= (axi_slave12)
`endif // ATCBMC300_SLV12_SUPPORT
`ifdef ATCBMC300_SLV13_SUPPORT
	.ds13_arvalid(ds13_arvalid), // (axi_monitor_s13,axi_slave13,bench) <= (bmc300)
	.ds13_arready(ds13_arready), // (axi_monitor_s13,bench,bmc300) <= (axi_slave13)
	.ds13_awvalid(ds13_awvalid), // (axi_monitor_s13,axi_slave13,bench) <= (bmc300)
	.ds13_awready(ds13_awready), // (axi_monitor_s13,bench,bmc300) <= (axi_slave13)
`endif // ATCBMC300_SLV13_SUPPORT
`ifdef ATCBMC300_SLV14_SUPPORT
	.ds14_arvalid(ds14_arvalid), // (axi_monitor_s14,axi_slave14,bench) <= (bmc300)
	.ds14_arready(ds14_arready), // (axi_monitor_s14,bench,bmc300) <= (axi_slave14)
	.ds14_awvalid(ds14_awvalid), // (axi_monitor_s14,axi_slave14,bench) <= (bmc300)
	.ds14_awready(ds14_awready), // (axi_monitor_s14,bench,bmc300) <= (axi_slave14)
`endif // ATCBMC300_SLV14_SUPPORT
`ifdef ATCBMC300_SLV15_SUPPORT
	.ds15_arvalid(ds15_arvalid), // (axi_monitor_s15,axi_slave15,bench) <= (bmc300)
	.ds15_arready(ds15_arready), // (axi_monitor_s15,bench,bmc300) <= (axi_slave15)
	.ds15_awvalid(ds15_awvalid), // (axi_monitor_s15,axi_slave15,bench) <= (bmc300)
	.ds15_awready(ds15_awready), // (axi_monitor_s15,bench,bmc300) <= (axi_slave15)
`endif // ATCBMC300_SLV15_SUPPORT
`ifdef ATCBMC300_SLV16_SUPPORT
	.ds16_arvalid(ds16_arvalid), // (axi_monitor_s16,axi_slave16,bench) <= (bmc300)
	.ds16_arready(ds16_arready), // (axi_monitor_s16,bench,bmc300) <= (axi_slave16)
	.ds16_awvalid(ds16_awvalid), // (axi_monitor_s16,axi_slave16,bench) <= (bmc300)
	.ds16_awready(ds16_awready), // (axi_monitor_s16,bench,bmc300) <= (axi_slave16)
`endif // ATCBMC300_SLV16_SUPPORT
`ifdef ATCBMC300_SLV17_SUPPORT
	.ds17_arvalid(ds17_arvalid), // (axi_monitor_s17,axi_slave17,bench) <= (bmc300)
	.ds17_arready(ds17_arready), // (axi_monitor_s17,bench,bmc300) <= (axi_slave17)
	.ds17_awvalid(ds17_awvalid), // (axi_monitor_s17,axi_slave17,bench) <= (bmc300)
	.ds17_awready(ds17_awready), // (axi_monitor_s17,bench,bmc300) <= (axi_slave17)
`endif // ATCBMC300_SLV17_SUPPORT
`ifdef ATCBMC300_SLV18_SUPPORT
	.ds18_arvalid(ds18_arvalid), // (axi_monitor_s18,axi_slave18,bench) <= (bmc300)
	.ds18_arready(ds18_arready), // (axi_monitor_s18,bench,bmc300) <= (axi_slave18)
	.ds18_awvalid(ds18_awvalid), // (axi_monitor_s18,axi_slave18,bench) <= (bmc300)
	.ds18_awready(ds18_awready), // (axi_monitor_s18,bench,bmc300) <= (axi_slave18)
`endif // ATCBMC300_SLV18_SUPPORT
`ifdef ATCBMC300_SLV19_SUPPORT
	.ds19_arvalid(ds19_arvalid), // (axi_monitor_s19,axi_slave19,bench) <= (bmc300)
	.ds19_arready(ds19_arready), // (axi_monitor_s19,bench,bmc300) <= (axi_slave19)
	.ds19_awvalid(ds19_awvalid), // (axi_monitor_s19,axi_slave19,bench) <= (bmc300)
	.ds19_awready(ds19_awready), // (axi_monitor_s19,bench,bmc300) <= (axi_slave19)
`endif // ATCBMC300_SLV19_SUPPORT
`ifdef ATCBMC300_SLV20_SUPPORT
	.ds20_arvalid(ds20_arvalid), // (axi_monitor_s20,axi_slave20,bench) <= (bmc300)
	.ds20_arready(ds20_arready), // (axi_monitor_s20,bench,bmc300) <= (axi_slave20)
	.ds20_awvalid(ds20_awvalid), // (axi_monitor_s20,axi_slave20,bench) <= (bmc300)
	.ds20_awready(ds20_awready), // (axi_monitor_s20,bench,bmc300) <= (axi_slave20)
`endif // ATCBMC300_SLV20_SUPPORT
`ifdef ATCBMC300_SLV21_SUPPORT
	.ds21_arvalid(ds21_arvalid), // (axi_monitor_s21,axi_slave21,bench) <= (bmc300)
	.ds21_arready(ds21_arready), // (axi_monitor_s21,bench,bmc300) <= (axi_slave21)
	.ds21_awvalid(ds21_awvalid), // (axi_monitor_s21,axi_slave21,bench) <= (bmc300)
	.ds21_awready(ds21_awready), // (axi_monitor_s21,bench,bmc300) <= (axi_slave21)
`endif // ATCBMC300_SLV21_SUPPORT
`ifdef ATCBMC300_SLV22_SUPPORT
	.ds22_arvalid(ds22_arvalid), // (axi_monitor_s22,axi_slave22,bench) <= (bmc300)
	.ds22_arready(ds22_arready), // (axi_monitor_s22,bench,bmc300) <= (axi_slave22)
	.ds22_awvalid(ds22_awvalid), // (axi_monitor_s22,axi_slave22,bench) <= (bmc300)
	.ds22_awready(ds22_awready), // (axi_monitor_s22,bench,bmc300) <= (axi_slave22)
`endif // ATCBMC300_SLV22_SUPPORT
`ifdef ATCBMC300_SLV23_SUPPORT
	.ds23_arvalid(ds23_arvalid), // (axi_monitor_s23,axi_slave23,bench) <= (bmc300)
	.ds23_arready(ds23_arready), // (axi_monitor_s23,bench,bmc300) <= (axi_slave23)
	.ds23_awvalid(ds23_awvalid), // (axi_monitor_s23,axi_slave23,bench) <= (bmc300)
	.ds23_awready(ds23_awready), // (axi_monitor_s23,bench,bmc300) <= (axi_slave23)
`endif // ATCBMC300_SLV23_SUPPORT
`ifdef ATCBMC300_SLV24_SUPPORT
	.ds24_arvalid(ds24_arvalid), // (axi_monitor_s24,axi_slave24,bench) <= (bmc300)
	.ds24_arready(ds24_arready), // (axi_monitor_s24,bench,bmc300) <= (axi_slave24)
	.ds24_awvalid(ds24_awvalid), // (axi_monitor_s24,axi_slave24,bench) <= (bmc300)
	.ds24_awready(ds24_awready), // (axi_monitor_s24,bench,bmc300) <= (axi_slave24)
`endif // ATCBMC300_SLV24_SUPPORT
`ifdef ATCBMC300_SLV25_SUPPORT
	.ds25_arvalid(ds25_arvalid), // (axi_monitor_s25,axi_slave25,bench) <= (bmc300)
	.ds25_arready(ds25_arready), // (axi_monitor_s25,bench,bmc300) <= (axi_slave25)
	.ds25_awvalid(ds25_awvalid), // (axi_monitor_s25,axi_slave25,bench) <= (bmc300)
	.ds25_awready(ds25_awready), // (axi_monitor_s25,bench,bmc300) <= (axi_slave25)
`endif // ATCBMC300_SLV25_SUPPORT
`ifdef ATCBMC300_SLV26_SUPPORT
	.ds26_arvalid(ds26_arvalid), // (axi_monitor_s26,axi_slave26,bench) <= (bmc300)
	.ds26_arready(ds26_arready), // (axi_monitor_s26,bench,bmc300) <= (axi_slave26)
	.ds26_awvalid(ds26_awvalid), // (axi_monitor_s26,axi_slave26,bench) <= (bmc300)
	.ds26_awready(ds26_awready), // (axi_monitor_s26,bench,bmc300) <= (axi_slave26)
`endif // ATCBMC300_SLV26_SUPPORT
`ifdef ATCBMC300_SLV27_SUPPORT
	.ds27_arvalid(ds27_arvalid), // (axi_monitor_s27,axi_slave27,bench) <= (bmc300)
	.ds27_arready(ds27_arready), // (axi_monitor_s27,bench,bmc300) <= (axi_slave27)
	.ds27_awvalid(ds27_awvalid), // (axi_monitor_s27,axi_slave27,bench) <= (bmc300)
	.ds27_awready(ds27_awready), // (axi_monitor_s27,bench,bmc300) <= (axi_slave27)
`endif // ATCBMC300_SLV27_SUPPORT
`ifdef ATCBMC300_SLV28_SUPPORT
	.ds28_arvalid(ds28_arvalid), // (axi_monitor_s28,axi_slave28,bench) <= (bmc300)
	.ds28_arready(ds28_arready), // (axi_monitor_s28,bench,bmc300) <= (axi_slave28)
	.ds28_awvalid(ds28_awvalid), // (axi_monitor_s28,axi_slave28,bench) <= (bmc300)
	.ds28_awready(ds28_awready), // (axi_monitor_s28,bench,bmc300) <= (axi_slave28)
`endif // ATCBMC300_SLV28_SUPPORT
`ifdef ATCBMC300_SLV29_SUPPORT
	.ds29_arvalid(ds29_arvalid), // (axi_monitor_s29,axi_slave29,bench) <= (bmc300)
	.ds29_arready(ds29_arready), // (axi_monitor_s29,bench,bmc300) <= (axi_slave29)
	.ds29_awvalid(ds29_awvalid), // (axi_monitor_s29,axi_slave29,bench) <= (bmc300)
	.ds29_awready(ds29_awready), // (axi_monitor_s29,bench,bmc300) <= (axi_slave29)
`endif // ATCBMC300_SLV29_SUPPORT
`ifdef ATCBMC300_SLV30_SUPPORT
	.ds30_arvalid(ds30_arvalid), // (axi_monitor_s30,axi_slave30,bench) <= (bmc300)
	.ds30_arready(ds30_arready), // (axi_monitor_s30,bench,bmc300) <= (axi_slave30)
	.ds30_awvalid(ds30_awvalid), // (axi_monitor_s30,axi_slave30,bench) <= (bmc300)
	.ds30_awready(ds30_awready), // (axi_monitor_s30,bench,bmc300) <= (axi_slave30)
`endif // ATCBMC300_SLV30_SUPPORT
`ifdef ATCBMC300_SLV31_SUPPORT
	.ds31_arvalid(ds31_arvalid), // (axi_monitor_s31,axi_slave31,bench) <= (bmc300)
	.ds31_arready(ds31_arready), // (axi_monitor_s31,bench,bmc300) <= (axi_slave31)
	.ds31_awvalid(ds31_awvalid), // (axi_monitor_s31,axi_slave31,bench) <= (bmc300)
	.ds31_awready(ds31_awready), // (axi_monitor_s31,bench,bmc300) <= (axi_slave31)
`endif // ATCBMC300_SLV31_SUPPORT
	.aclk        (aclk        ), // (bench) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300)
	.aresetn     (aresetn     )  // (bench) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300)
); // end of bench

`ifdef ATCBMC300_MST0_SUPPORT
defparam axi_master0.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master0.ADDR_START = 0;
defparam axi_master0.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master0.AXI4 = 1'b1;
defparam axi_master0.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master0.DATA_WIDTH = DATA_SIZE;
defparam axi_master0.DELAY_MAX = `ifdef NDS_MST0_DELAY_MAX `NDS_MST0_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master0.ID_WIDTH = US_ID_WIDTH;
defparam axi_master0.MAX_BUF_DEPTH = 256;
defparam axi_master0.MODEL_ID = 0;
defparam axi_master0.TRANS_NUM = `ifdef NDS_MST0_TRANS_NUM `NDS_MST0_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master0.UNALIGN_SUPPORT = 1'b1;
defparam axi_master0.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master0 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us0_awid                  ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.awaddr  (us0_awaddr                ), // (axi_master0) => (axi_monitor_m0,bench,bmc300)
	.awlen   (us0_awlen                 ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.awsize  (us0_awsize                ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.awburst (us0_awburst               ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.awlock  ({us0_awlock_b1,us0_awlock}), // () => ()
	.awcache (us0_awcache               ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.awprot  (us0_awprot                ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.awvalid (us0_awvalid               ), // (axi_master0) => (axi_monitor_m0,bench,bmc300)
	.awready (us0_awready               ), // (axi_master0,axi_monitor_m0,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us0_wid                   ), // (axi_master0) => (axi_monitor_m0)
	.wdata   (us0_wdata                 ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.wstrb   (us0_wstrb                 ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.wlast   (us0_wlast                 ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.wvalid  (us0_wvalid                ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.wready  (us0_wready                ), // (axi_master0,axi_monitor_m0) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us0_bid                   ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.bresp   (us0_bresp                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.bvalid  (us0_bvalid                ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.bready  (us0_bready                ), // (axi_master0) => (axi_monitor_m0,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us0_arid                  ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.araddr  (us0_araddr                ), // (axi_master0) => (axi_monitor_m0,bench,bmc300)
	.arlen   (us0_arlen                 ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.arsize  (us0_arsize                ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.arburst (us0_arburst               ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.arlock  ({us0_arlock_b1,us0_arlock}), // () => ()
	.arcache (us0_arcache               ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.arprot  (us0_arprot                ), // (axi_master0) => (axi_monitor_m0,bmc300)
	.arvalid (us0_arvalid               ), // (axi_master0) => (axi_monitor_m0,bench,bmc300)
	.arready (us0_arready               ), // (axi_master0,axi_monitor_m0,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us0_rid                   ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rdata   (us0_rdata                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rresp   (us0_rresp                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rlast   (us0_rlast                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rvalid  (us0_rvalid                ), // (axi_master0,axi_monitor_m0) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us0_rready                )  // (axi_master0) => (axi_monitor_m0,bmc300)
); // end of axi_master0

defparam axi_monitor_m0.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m0.AXI4 = 1'b1;
defparam axi_monitor_m0.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m0.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m0.MASTER_ID = 0;
defparam axi_monitor_m0.SLAVE_ID = 0;
axi_monitor axi_monitor_m0 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us0_awid                  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.awaddr  (us0_awaddr                ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.awlen   (us0_awlen                 ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.awsize  (us0_awsize                ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.awburst (us0_awburst               ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.awlock  ({us0_awlock_b1,us0_awlock}), // () <= ()
	.awcache (us0_awcache               ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.awprot  (us0_awprot                ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.awvalid (us0_awvalid               ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.awready (us0_awready               ), // (axi_master0,axi_monitor_m0,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us0_wid                   ), // (axi_monitor_m0) <= (axi_master0)
	.wdata   (us0_wdata                 ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.wstrb   (us0_wstrb                 ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.wlast   (us0_wlast                 ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.wvalid  (us0_wvalid                ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.wready  (us0_wready                ), // (axi_master0,axi_monitor_m0) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us0_bid                   ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.bresp   (us0_bresp                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.bvalid  (us0_bvalid                ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.bready  (us0_bready                ), // (axi_monitor_m0,bmc300) <= (axi_master0)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us0_arid                  ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.araddr  (us0_araddr                ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.arlen   (us0_arlen                 ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.arsize  (us0_arsize                ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.arburst (us0_arburst               ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.arlock  ({us0_arlock_b1,us0_arlock}), // () <= ()
	.arcache (us0_arcache               ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.arprot  (us0_arprot                ), // (axi_monitor_m0,bmc300) <= (axi_master0)
	.arvalid (us0_arvalid               ), // (axi_monitor_m0,bench,bmc300) <= (axi_master0)
	.arready (us0_arready               ), // (axi_master0,axi_monitor_m0,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us0_rid                   ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rdata   (us0_rdata                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rresp   (us0_rresp                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rlast   (us0_rlast                 ), // (axi_master0,axi_monitor_m0) <= (bmc300)
	.rvalid  (us0_rvalid                ), // (axi_master0,axi_monitor_m0) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us0_rready                )  // (axi_monitor_m0,bmc300) <= (axi_master0)
); // end of axi_monitor_m0

`endif // ATCBMC300_MST0_SUPPORT
`ifdef ATCBMC300_MST1_SUPPORT
defparam axi_master1.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master1.ADDR_START = 0;
defparam axi_master1.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master1.AXI4 = 1'b1;
defparam axi_master1.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master1.DATA_WIDTH = DATA_SIZE;
defparam axi_master1.DELAY_MAX = `ifdef NDS_MST1_DELAY_MAX `NDS_MST1_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master1.ID_WIDTH = US_ID_WIDTH;
defparam axi_master1.MAX_BUF_DEPTH = 256;
defparam axi_master1.MODEL_ID = 1;
defparam axi_master1.TRANS_NUM = `ifdef NDS_MST1_TRANS_NUM `NDS_MST1_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master1.UNALIGN_SUPPORT = 1'b1;
defparam axi_master1.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master1 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us1_awid                  ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.awaddr  (us1_awaddr                ), // (axi_master1) => (axi_monitor_m1,bench,bmc300)
	.awlen   (us1_awlen                 ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.awsize  (us1_awsize                ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.awburst (us1_awburst               ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.awlock  ({us1_awlock_b1,us1_awlock}), // () => ()
	.awcache (us1_awcache               ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.awprot  (us1_awprot                ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.awvalid (us1_awvalid               ), // (axi_master1) => (axi_monitor_m1,bench,bmc300)
	.awready (us1_awready               ), // (axi_master1,axi_monitor_m1,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us1_wid                   ), // (axi_master1) => (axi_monitor_m1)
	.wdata   (us1_wdata                 ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.wstrb   (us1_wstrb                 ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.wlast   (us1_wlast                 ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.wvalid  (us1_wvalid                ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.wready  (us1_wready                ), // (axi_master1,axi_monitor_m1) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us1_bid                   ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.bresp   (us1_bresp                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.bvalid  (us1_bvalid                ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.bready  (us1_bready                ), // (axi_master1) => (axi_monitor_m1,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us1_arid                  ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.araddr  (us1_araddr                ), // (axi_master1) => (axi_monitor_m1,bench,bmc300)
	.arlen   (us1_arlen                 ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.arsize  (us1_arsize                ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.arburst (us1_arburst               ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.arlock  ({us1_arlock_b1,us1_arlock}), // () => ()
	.arcache (us1_arcache               ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.arprot  (us1_arprot                ), // (axi_master1) => (axi_monitor_m1,bmc300)
	.arvalid (us1_arvalid               ), // (axi_master1) => (axi_monitor_m1,bench,bmc300)
	.arready (us1_arready               ), // (axi_master1,axi_monitor_m1,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us1_rid                   ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rdata   (us1_rdata                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rresp   (us1_rresp                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rlast   (us1_rlast                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rvalid  (us1_rvalid                ), // (axi_master1,axi_monitor_m1) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us1_rready                )  // (axi_master1) => (axi_monitor_m1,bmc300)
); // end of axi_master1

defparam axi_monitor_m1.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m1.AXI4 = 1'b1;
defparam axi_monitor_m1.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m1.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m1.MASTER_ID = 1;
defparam axi_monitor_m1.SLAVE_ID = 1;
axi_monitor axi_monitor_m1 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us1_awid                  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.awaddr  (us1_awaddr                ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.awlen   (us1_awlen                 ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.awsize  (us1_awsize                ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.awburst (us1_awburst               ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.awlock  ({us1_awlock_b1,us1_awlock}), // () <= ()
	.awcache (us1_awcache               ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.awprot  (us1_awprot                ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.awvalid (us1_awvalid               ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.awready (us1_awready               ), // (axi_master1,axi_monitor_m1,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us1_wid                   ), // (axi_monitor_m1) <= (axi_master1)
	.wdata   (us1_wdata                 ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.wstrb   (us1_wstrb                 ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.wlast   (us1_wlast                 ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.wvalid  (us1_wvalid                ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.wready  (us1_wready                ), // (axi_master1,axi_monitor_m1) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us1_bid                   ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.bresp   (us1_bresp                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.bvalid  (us1_bvalid                ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.bready  (us1_bready                ), // (axi_monitor_m1,bmc300) <= (axi_master1)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us1_arid                  ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.araddr  (us1_araddr                ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.arlen   (us1_arlen                 ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.arsize  (us1_arsize                ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.arburst (us1_arburst               ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.arlock  ({us1_arlock_b1,us1_arlock}), // () <= ()
	.arcache (us1_arcache               ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.arprot  (us1_arprot                ), // (axi_monitor_m1,bmc300) <= (axi_master1)
	.arvalid (us1_arvalid               ), // (axi_monitor_m1,bench,bmc300) <= (axi_master1)
	.arready (us1_arready               ), // (axi_master1,axi_monitor_m1,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us1_rid                   ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rdata   (us1_rdata                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rresp   (us1_rresp                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rlast   (us1_rlast                 ), // (axi_master1,axi_monitor_m1) <= (bmc300)
	.rvalid  (us1_rvalid                ), // (axi_master1,axi_monitor_m1) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us1_rready                )  // (axi_monitor_m1,bmc300) <= (axi_master1)
); // end of axi_monitor_m1

`endif // ATCBMC300_MST1_SUPPORT
`ifdef ATCBMC300_MST2_SUPPORT
defparam axi_master2.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master2.ADDR_START = 0;
defparam axi_master2.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master2.AXI4 = 1'b1;
defparam axi_master2.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master2.DATA_WIDTH = DATA_SIZE;
defparam axi_master2.DELAY_MAX = `ifdef NDS_MST2_DELAY_MAX `NDS_MST2_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master2.ID_WIDTH = US_ID_WIDTH;
defparam axi_master2.MAX_BUF_DEPTH = 256;
defparam axi_master2.MODEL_ID = 2;
defparam axi_master2.TRANS_NUM = `ifdef NDS_MST2_TRANS_NUM `NDS_MST2_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master2.UNALIGN_SUPPORT = 1'b1;
defparam axi_master2.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master2 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us2_awid                  ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.awaddr  (us2_awaddr                ), // (axi_master2) => (axi_monitor_m2,bench,bmc300)
	.awlen   (us2_awlen                 ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.awsize  (us2_awsize                ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.awburst (us2_awburst               ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.awlock  ({us2_awlock_b1,us2_awlock}), // () => ()
	.awcache (us2_awcache               ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.awprot  (us2_awprot                ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.awvalid (us2_awvalid               ), // (axi_master2) => (axi_monitor_m2,bench,bmc300)
	.awready (us2_awready               ), // (axi_master2,axi_monitor_m2,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us2_wid                   ), // (axi_master2) => (axi_monitor_m2)
	.wdata   (us2_wdata                 ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.wstrb   (us2_wstrb                 ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.wlast   (us2_wlast                 ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.wvalid  (us2_wvalid                ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.wready  (us2_wready                ), // (axi_master2,axi_monitor_m2) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us2_bid                   ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.bresp   (us2_bresp                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.bvalid  (us2_bvalid                ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.bready  (us2_bready                ), // (axi_master2) => (axi_monitor_m2,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us2_arid                  ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.araddr  (us2_araddr                ), // (axi_master2) => (axi_monitor_m2,bench,bmc300)
	.arlen   (us2_arlen                 ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.arsize  (us2_arsize                ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.arburst (us2_arburst               ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.arlock  ({us2_arlock_b1,us2_arlock}), // () => ()
	.arcache (us2_arcache               ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.arprot  (us2_arprot                ), // (axi_master2) => (axi_monitor_m2,bmc300)
	.arvalid (us2_arvalid               ), // (axi_master2) => (axi_monitor_m2,bench,bmc300)
	.arready (us2_arready               ), // (axi_master2,axi_monitor_m2,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us2_rid                   ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rdata   (us2_rdata                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rresp   (us2_rresp                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rlast   (us2_rlast                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rvalid  (us2_rvalid                ), // (axi_master2,axi_monitor_m2) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us2_rready                )  // (axi_master2) => (axi_monitor_m2,bmc300)
); // end of axi_master2

defparam axi_monitor_m2.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m2.AXI4 = 1'b1;
defparam axi_monitor_m2.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m2.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m2.MASTER_ID = 2;
defparam axi_monitor_m2.SLAVE_ID = 2;
axi_monitor axi_monitor_m2 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us2_awid                  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.awaddr  (us2_awaddr                ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.awlen   (us2_awlen                 ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.awsize  (us2_awsize                ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.awburst (us2_awburst               ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.awlock  ({us2_awlock_b1,us2_awlock}), // () <= ()
	.awcache (us2_awcache               ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.awprot  (us2_awprot                ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.awvalid (us2_awvalid               ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.awready (us2_awready               ), // (axi_master2,axi_monitor_m2,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us2_wid                   ), // (axi_monitor_m2) <= (axi_master2)
	.wdata   (us2_wdata                 ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.wstrb   (us2_wstrb                 ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.wlast   (us2_wlast                 ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.wvalid  (us2_wvalid                ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.wready  (us2_wready                ), // (axi_master2,axi_monitor_m2) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us2_bid                   ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.bresp   (us2_bresp                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.bvalid  (us2_bvalid                ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.bready  (us2_bready                ), // (axi_monitor_m2,bmc300) <= (axi_master2)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us2_arid                  ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.araddr  (us2_araddr                ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.arlen   (us2_arlen                 ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.arsize  (us2_arsize                ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.arburst (us2_arburst               ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.arlock  ({us2_arlock_b1,us2_arlock}), // () <= ()
	.arcache (us2_arcache               ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.arprot  (us2_arprot                ), // (axi_monitor_m2,bmc300) <= (axi_master2)
	.arvalid (us2_arvalid               ), // (axi_monitor_m2,bench,bmc300) <= (axi_master2)
	.arready (us2_arready               ), // (axi_master2,axi_monitor_m2,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us2_rid                   ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rdata   (us2_rdata                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rresp   (us2_rresp                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rlast   (us2_rlast                 ), // (axi_master2,axi_monitor_m2) <= (bmc300)
	.rvalid  (us2_rvalid                ), // (axi_master2,axi_monitor_m2) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us2_rready                )  // (axi_monitor_m2,bmc300) <= (axi_master2)
); // end of axi_monitor_m2

`endif // ATCBMC300_MST2_SUPPORT
`ifdef ATCBMC300_MST3_SUPPORT
defparam axi_master3.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master3.ADDR_START = 0;
defparam axi_master3.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master3.AXI4 = 1'b1;
defparam axi_master3.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master3.DATA_WIDTH = DATA_SIZE;
defparam axi_master3.DELAY_MAX = `ifdef NDS_MST3_DELAY_MAX `NDS_MST3_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master3.ID_WIDTH = US_ID_WIDTH;
defparam axi_master3.MAX_BUF_DEPTH = 256;
defparam axi_master3.MODEL_ID = 3;
defparam axi_master3.TRANS_NUM = `ifdef NDS_MST3_TRANS_NUM `NDS_MST3_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master3.UNALIGN_SUPPORT = 1'b1;
defparam axi_master3.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master3 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us3_awid                  ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.awaddr  (us3_awaddr                ), // (axi_master3) => (axi_monitor_m3,bench,bmc300)
	.awlen   (us3_awlen                 ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.awsize  (us3_awsize                ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.awburst (us3_awburst               ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.awlock  ({us3_awlock_b1,us3_awlock}), // () => ()
	.awcache (us3_awcache               ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.awprot  (us3_awprot                ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.awvalid (us3_awvalid               ), // (axi_master3) => (axi_monitor_m3,bench,bmc300)
	.awready (us3_awready               ), // (axi_master3,axi_monitor_m3,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us3_wid                   ), // (axi_master3) => (axi_monitor_m3)
	.wdata   (us3_wdata                 ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.wstrb   (us3_wstrb                 ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.wlast   (us3_wlast                 ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.wvalid  (us3_wvalid                ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.wready  (us3_wready                ), // (axi_master3,axi_monitor_m3) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us3_bid                   ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.bresp   (us3_bresp                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.bvalid  (us3_bvalid                ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.bready  (us3_bready                ), // (axi_master3) => (axi_monitor_m3,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us3_arid                  ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.araddr  (us3_araddr                ), // (axi_master3) => (axi_monitor_m3,bench,bmc300)
	.arlen   (us3_arlen                 ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.arsize  (us3_arsize                ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.arburst (us3_arburst               ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.arlock  ({us3_arlock_b1,us3_arlock}), // () => ()
	.arcache (us3_arcache               ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.arprot  (us3_arprot                ), // (axi_master3) => (axi_monitor_m3,bmc300)
	.arvalid (us3_arvalid               ), // (axi_master3) => (axi_monitor_m3,bench,bmc300)
	.arready (us3_arready               ), // (axi_master3,axi_monitor_m3,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us3_rid                   ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rdata   (us3_rdata                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rresp   (us3_rresp                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rlast   (us3_rlast                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rvalid  (us3_rvalid                ), // (axi_master3,axi_monitor_m3) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us3_rready                )  // (axi_master3) => (axi_monitor_m3,bmc300)
); // end of axi_master3

defparam axi_monitor_m3.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m3.AXI4 = 1'b1;
defparam axi_monitor_m3.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m3.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m3.MASTER_ID = 3;
defparam axi_monitor_m3.SLAVE_ID = 3;
axi_monitor axi_monitor_m3 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us3_awid                  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.awaddr  (us3_awaddr                ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.awlen   (us3_awlen                 ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.awsize  (us3_awsize                ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.awburst (us3_awburst               ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.awlock  ({us3_awlock_b1,us3_awlock}), // () <= ()
	.awcache (us3_awcache               ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.awprot  (us3_awprot                ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.awvalid (us3_awvalid               ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.awready (us3_awready               ), // (axi_master3,axi_monitor_m3,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us3_wid                   ), // (axi_monitor_m3) <= (axi_master3)
	.wdata   (us3_wdata                 ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.wstrb   (us3_wstrb                 ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.wlast   (us3_wlast                 ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.wvalid  (us3_wvalid                ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.wready  (us3_wready                ), // (axi_master3,axi_monitor_m3) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us3_bid                   ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.bresp   (us3_bresp                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.bvalid  (us3_bvalid                ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.bready  (us3_bready                ), // (axi_monitor_m3,bmc300) <= (axi_master3)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us3_arid                  ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.araddr  (us3_araddr                ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.arlen   (us3_arlen                 ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.arsize  (us3_arsize                ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.arburst (us3_arburst               ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.arlock  ({us3_arlock_b1,us3_arlock}), // () <= ()
	.arcache (us3_arcache               ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.arprot  (us3_arprot                ), // (axi_monitor_m3,bmc300) <= (axi_master3)
	.arvalid (us3_arvalid               ), // (axi_monitor_m3,bench,bmc300) <= (axi_master3)
	.arready (us3_arready               ), // (axi_master3,axi_monitor_m3,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us3_rid                   ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rdata   (us3_rdata                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rresp   (us3_rresp                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rlast   (us3_rlast                 ), // (axi_master3,axi_monitor_m3) <= (bmc300)
	.rvalid  (us3_rvalid                ), // (axi_master3,axi_monitor_m3) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us3_rready                )  // (axi_monitor_m3,bmc300) <= (axi_master3)
); // end of axi_monitor_m3

`endif // ATCBMC300_MST3_SUPPORT
`ifdef ATCBMC300_MST4_SUPPORT
defparam axi_master4.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master4.ADDR_START = 0;
defparam axi_master4.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master4.AXI4 = 1'b1;
defparam axi_master4.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master4.DATA_WIDTH = DATA_SIZE;
defparam axi_master4.DELAY_MAX = `ifdef NDS_MST4_DELAY_MAX `NDS_MST4_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master4.ID_WIDTH = US_ID_WIDTH;
defparam axi_master4.MAX_BUF_DEPTH = 256;
defparam axi_master4.MODEL_ID = 4;
defparam axi_master4.TRANS_NUM = `ifdef NDS_MST4_TRANS_NUM `NDS_MST4_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master4.UNALIGN_SUPPORT = 1'b1;
defparam axi_master4.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master4 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us4_awid                  ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.awaddr  (us4_awaddr                ), // (axi_master4) => (axi_monitor_m4,bench,bmc300)
	.awlen   (us4_awlen                 ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.awsize  (us4_awsize                ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.awburst (us4_awburst               ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.awlock  ({us4_awlock_b1,us4_awlock}), // () => ()
	.awcache (us4_awcache               ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.awprot  (us4_awprot                ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.awvalid (us4_awvalid               ), // (axi_master4) => (axi_monitor_m4,bench,bmc300)
	.awready (us4_awready               ), // (axi_master4,axi_monitor_m4,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us4_wid                   ), // (axi_master4) => (axi_monitor_m4)
	.wdata   (us4_wdata                 ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.wstrb   (us4_wstrb                 ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.wlast   (us4_wlast                 ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.wvalid  (us4_wvalid                ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.wready  (us4_wready                ), // (axi_master4,axi_monitor_m4) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us4_bid                   ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.bresp   (us4_bresp                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.bvalid  (us4_bvalid                ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.bready  (us4_bready                ), // (axi_master4) => (axi_monitor_m4,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us4_arid                  ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.araddr  (us4_araddr                ), // (axi_master4) => (axi_monitor_m4,bench,bmc300)
	.arlen   (us4_arlen                 ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.arsize  (us4_arsize                ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.arburst (us4_arburst               ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.arlock  ({us4_arlock_b1,us4_arlock}), // () => ()
	.arcache (us4_arcache               ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.arprot  (us4_arprot                ), // (axi_master4) => (axi_monitor_m4,bmc300)
	.arvalid (us4_arvalid               ), // (axi_master4) => (axi_monitor_m4,bench,bmc300)
	.arready (us4_arready               ), // (axi_master4,axi_monitor_m4,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us4_rid                   ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rdata   (us4_rdata                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rresp   (us4_rresp                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rlast   (us4_rlast                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rvalid  (us4_rvalid                ), // (axi_master4,axi_monitor_m4) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us4_rready                )  // (axi_master4) => (axi_monitor_m4,bmc300)
); // end of axi_master4

defparam axi_monitor_m4.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m4.AXI4 = 1'b1;
defparam axi_monitor_m4.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m4.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m4.MASTER_ID = 4;
defparam axi_monitor_m4.SLAVE_ID = 4;
axi_monitor axi_monitor_m4 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us4_awid                  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.awaddr  (us4_awaddr                ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.awlen   (us4_awlen                 ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.awsize  (us4_awsize                ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.awburst (us4_awburst               ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.awlock  ({us4_awlock_b1,us4_awlock}), // () <= ()
	.awcache (us4_awcache               ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.awprot  (us4_awprot                ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.awvalid (us4_awvalid               ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.awready (us4_awready               ), // (axi_master4,axi_monitor_m4,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us4_wid                   ), // (axi_monitor_m4) <= (axi_master4)
	.wdata   (us4_wdata                 ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.wstrb   (us4_wstrb                 ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.wlast   (us4_wlast                 ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.wvalid  (us4_wvalid                ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.wready  (us4_wready                ), // (axi_master4,axi_monitor_m4) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us4_bid                   ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.bresp   (us4_bresp                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.bvalid  (us4_bvalid                ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.bready  (us4_bready                ), // (axi_monitor_m4,bmc300) <= (axi_master4)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us4_arid                  ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.araddr  (us4_araddr                ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.arlen   (us4_arlen                 ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.arsize  (us4_arsize                ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.arburst (us4_arburst               ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.arlock  ({us4_arlock_b1,us4_arlock}), // () <= ()
	.arcache (us4_arcache               ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.arprot  (us4_arprot                ), // (axi_monitor_m4,bmc300) <= (axi_master4)
	.arvalid (us4_arvalid               ), // (axi_monitor_m4,bench,bmc300) <= (axi_master4)
	.arready (us4_arready               ), // (axi_master4,axi_monitor_m4,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us4_rid                   ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rdata   (us4_rdata                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rresp   (us4_rresp                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rlast   (us4_rlast                 ), // (axi_master4,axi_monitor_m4) <= (bmc300)
	.rvalid  (us4_rvalid                ), // (axi_master4,axi_monitor_m4) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us4_rready                )  // (axi_monitor_m4,bmc300) <= (axi_master4)
); // end of axi_monitor_m4

`endif // ATCBMC300_MST4_SUPPORT
`ifdef ATCBMC300_MST5_SUPPORT
defparam axi_master5.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master5.ADDR_START = 0;
defparam axi_master5.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master5.AXI4 = 1'b1;
defparam axi_master5.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master5.DATA_WIDTH = DATA_SIZE;
defparam axi_master5.DELAY_MAX = `ifdef NDS_MST5_DELAY_MAX `NDS_MST5_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master5.ID_WIDTH = US_ID_WIDTH;
defparam axi_master5.MAX_BUF_DEPTH = 256;
defparam axi_master5.MODEL_ID = 5;
defparam axi_master5.TRANS_NUM = `ifdef NDS_MST5_TRANS_NUM `NDS_MST5_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master5.UNALIGN_SUPPORT = 1'b1;
defparam axi_master5.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master5 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us5_awid                  ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.awaddr  (us5_awaddr                ), // (axi_master5) => (axi_monitor_m5,bench,bmc300)
	.awlen   (us5_awlen                 ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.awsize  (us5_awsize                ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.awburst (us5_awburst               ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.awlock  ({us5_awlock_b1,us5_awlock}), // () => ()
	.awcache (us5_awcache               ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.awprot  (us5_awprot                ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.awvalid (us5_awvalid               ), // (axi_master5) => (axi_monitor_m5,bench,bmc300)
	.awready (us5_awready               ), // (axi_master5,axi_monitor_m5,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us5_wid                   ), // (axi_master5) => (axi_monitor_m5)
	.wdata   (us5_wdata                 ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.wstrb   (us5_wstrb                 ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.wlast   (us5_wlast                 ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.wvalid  (us5_wvalid                ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.wready  (us5_wready                ), // (axi_master5,axi_monitor_m5) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us5_bid                   ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.bresp   (us5_bresp                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.bvalid  (us5_bvalid                ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.bready  (us5_bready                ), // (axi_master5) => (axi_monitor_m5,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us5_arid                  ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.araddr  (us5_araddr                ), // (axi_master5) => (axi_monitor_m5,bench,bmc300)
	.arlen   (us5_arlen                 ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.arsize  (us5_arsize                ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.arburst (us5_arburst               ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.arlock  ({us5_arlock_b1,us5_arlock}), // () => ()
	.arcache (us5_arcache               ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.arprot  (us5_arprot                ), // (axi_master5) => (axi_monitor_m5,bmc300)
	.arvalid (us5_arvalid               ), // (axi_master5) => (axi_monitor_m5,bench,bmc300)
	.arready (us5_arready               ), // (axi_master5,axi_monitor_m5,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us5_rid                   ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rdata   (us5_rdata                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rresp   (us5_rresp                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rlast   (us5_rlast                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rvalid  (us5_rvalid                ), // (axi_master5,axi_monitor_m5) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us5_rready                )  // (axi_master5) => (axi_monitor_m5,bmc300)
); // end of axi_master5

defparam axi_monitor_m5.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m5.AXI4 = 1'b1;
defparam axi_monitor_m5.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m5.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m5.MASTER_ID = 5;
defparam axi_monitor_m5.SLAVE_ID = 5;
axi_monitor axi_monitor_m5 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us5_awid                  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.awaddr  (us5_awaddr                ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.awlen   (us5_awlen                 ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.awsize  (us5_awsize                ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.awburst (us5_awburst               ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.awlock  ({us5_awlock_b1,us5_awlock}), // () <= ()
	.awcache (us5_awcache               ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.awprot  (us5_awprot                ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.awvalid (us5_awvalid               ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.awready (us5_awready               ), // (axi_master5,axi_monitor_m5,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us5_wid                   ), // (axi_monitor_m5) <= (axi_master5)
	.wdata   (us5_wdata                 ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.wstrb   (us5_wstrb                 ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.wlast   (us5_wlast                 ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.wvalid  (us5_wvalid                ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.wready  (us5_wready                ), // (axi_master5,axi_monitor_m5) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us5_bid                   ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.bresp   (us5_bresp                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.bvalid  (us5_bvalid                ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.bready  (us5_bready                ), // (axi_monitor_m5,bmc300) <= (axi_master5)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us5_arid                  ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.araddr  (us5_araddr                ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.arlen   (us5_arlen                 ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.arsize  (us5_arsize                ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.arburst (us5_arburst               ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.arlock  ({us5_arlock_b1,us5_arlock}), // () <= ()
	.arcache (us5_arcache               ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.arprot  (us5_arprot                ), // (axi_monitor_m5,bmc300) <= (axi_master5)
	.arvalid (us5_arvalid               ), // (axi_monitor_m5,bench,bmc300) <= (axi_master5)
	.arready (us5_arready               ), // (axi_master5,axi_monitor_m5,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us5_rid                   ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rdata   (us5_rdata                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rresp   (us5_rresp                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rlast   (us5_rlast                 ), // (axi_master5,axi_monitor_m5) <= (bmc300)
	.rvalid  (us5_rvalid                ), // (axi_master5,axi_monitor_m5) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us5_rready                )  // (axi_monitor_m5,bmc300) <= (axi_master5)
); // end of axi_monitor_m5

`endif // ATCBMC300_MST5_SUPPORT
`ifdef ATCBMC300_MST6_SUPPORT
defparam axi_master6.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master6.ADDR_START = 0;
defparam axi_master6.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master6.AXI4 = 1'b1;
defparam axi_master6.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master6.DATA_WIDTH = DATA_SIZE;
defparam axi_master6.DELAY_MAX = `ifdef NDS_MST6_DELAY_MAX `NDS_MST6_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master6.ID_WIDTH = US_ID_WIDTH;
defparam axi_master6.MAX_BUF_DEPTH = 256;
defparam axi_master6.MODEL_ID = 6;
defparam axi_master6.TRANS_NUM = `ifdef NDS_MST6_TRANS_NUM `NDS_MST6_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master6.UNALIGN_SUPPORT = 1'b1;
defparam axi_master6.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master6 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us6_awid                  ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.awaddr  (us6_awaddr                ), // (axi_master6) => (axi_monitor_m6,bench,bmc300)
	.awlen   (us6_awlen                 ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.awsize  (us6_awsize                ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.awburst (us6_awburst               ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.awlock  ({us6_awlock_b1,us6_awlock}), // () => ()
	.awcache (us6_awcache               ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.awprot  (us6_awprot                ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.awvalid (us6_awvalid               ), // (axi_master6) => (axi_monitor_m6,bench,bmc300)
	.awready (us6_awready               ), // (axi_master6,axi_monitor_m6,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us6_wid                   ), // (axi_master6) => (axi_monitor_m6)
	.wdata   (us6_wdata                 ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.wstrb   (us6_wstrb                 ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.wlast   (us6_wlast                 ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.wvalid  (us6_wvalid                ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.wready  (us6_wready                ), // (axi_master6,axi_monitor_m6) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us6_bid                   ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.bresp   (us6_bresp                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.bvalid  (us6_bvalid                ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.bready  (us6_bready                ), // (axi_master6) => (axi_monitor_m6,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us6_arid                  ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.araddr  (us6_araddr                ), // (axi_master6) => (axi_monitor_m6,bench,bmc300)
	.arlen   (us6_arlen                 ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.arsize  (us6_arsize                ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.arburst (us6_arburst               ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.arlock  ({us6_arlock_b1,us6_arlock}), // () => ()
	.arcache (us6_arcache               ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.arprot  (us6_arprot                ), // (axi_master6) => (axi_monitor_m6,bmc300)
	.arvalid (us6_arvalid               ), // (axi_master6) => (axi_monitor_m6,bench,bmc300)
	.arready (us6_arready               ), // (axi_master6,axi_monitor_m6,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us6_rid                   ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rdata   (us6_rdata                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rresp   (us6_rresp                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rlast   (us6_rlast                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rvalid  (us6_rvalid                ), // (axi_master6,axi_monitor_m6) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us6_rready                )  // (axi_master6) => (axi_monitor_m6,bmc300)
); // end of axi_master6

defparam axi_monitor_m6.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m6.AXI4 = 1'b1;
defparam axi_monitor_m6.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m6.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m6.MASTER_ID = 6;
defparam axi_monitor_m6.SLAVE_ID = 6;
axi_monitor axi_monitor_m6 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us6_awid                  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.awaddr  (us6_awaddr                ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.awlen   (us6_awlen                 ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.awsize  (us6_awsize                ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.awburst (us6_awburst               ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.awlock  ({us6_awlock_b1,us6_awlock}), // () <= ()
	.awcache (us6_awcache               ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.awprot  (us6_awprot                ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.awvalid (us6_awvalid               ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.awready (us6_awready               ), // (axi_master6,axi_monitor_m6,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us6_wid                   ), // (axi_monitor_m6) <= (axi_master6)
	.wdata   (us6_wdata                 ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.wstrb   (us6_wstrb                 ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.wlast   (us6_wlast                 ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.wvalid  (us6_wvalid                ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.wready  (us6_wready                ), // (axi_master6,axi_monitor_m6) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us6_bid                   ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.bresp   (us6_bresp                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.bvalid  (us6_bvalid                ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.bready  (us6_bready                ), // (axi_monitor_m6,bmc300) <= (axi_master6)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us6_arid                  ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.araddr  (us6_araddr                ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.arlen   (us6_arlen                 ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.arsize  (us6_arsize                ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.arburst (us6_arburst               ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.arlock  ({us6_arlock_b1,us6_arlock}), // () <= ()
	.arcache (us6_arcache               ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.arprot  (us6_arprot                ), // (axi_monitor_m6,bmc300) <= (axi_master6)
	.arvalid (us6_arvalid               ), // (axi_monitor_m6,bench,bmc300) <= (axi_master6)
	.arready (us6_arready               ), // (axi_master6,axi_monitor_m6,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us6_rid                   ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rdata   (us6_rdata                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rresp   (us6_rresp                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rlast   (us6_rlast                 ), // (axi_master6,axi_monitor_m6) <= (bmc300)
	.rvalid  (us6_rvalid                ), // (axi_master6,axi_monitor_m6) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us6_rready                )  // (axi_monitor_m6,bmc300) <= (axi_master6)
); // end of axi_monitor_m6

`endif // ATCBMC300_MST6_SUPPORT
`ifdef ATCBMC300_MST7_SUPPORT
defparam axi_master7.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master7.ADDR_START = 0;
defparam axi_master7.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master7.AXI4 = 1'b1;
defparam axi_master7.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master7.DATA_WIDTH = DATA_SIZE;
defparam axi_master7.DELAY_MAX = `ifdef NDS_MST7_DELAY_MAX `NDS_MST7_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master7.ID_WIDTH = US_ID_WIDTH;
defparam axi_master7.MAX_BUF_DEPTH = 256;
defparam axi_master7.MODEL_ID = 7;
defparam axi_master7.TRANS_NUM = `ifdef NDS_MST7_TRANS_NUM `NDS_MST7_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master7.UNALIGN_SUPPORT = 1'b1;
defparam axi_master7.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master7 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us7_awid                  ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.awaddr  (us7_awaddr                ), // (axi_master7) => (axi_monitor_m7,bench,bmc300)
	.awlen   (us7_awlen                 ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.awsize  (us7_awsize                ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.awburst (us7_awburst               ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.awlock  ({us7_awlock_b1,us7_awlock}), // () => ()
	.awcache (us7_awcache               ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.awprot  (us7_awprot                ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.awvalid (us7_awvalid               ), // (axi_master7) => (axi_monitor_m7,bench,bmc300)
	.awready (us7_awready               ), // (axi_master7,axi_monitor_m7,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us7_wid                   ), // (axi_master7) => (axi_monitor_m7)
	.wdata   (us7_wdata                 ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.wstrb   (us7_wstrb                 ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.wlast   (us7_wlast                 ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.wvalid  (us7_wvalid                ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.wready  (us7_wready                ), // (axi_master7,axi_monitor_m7) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us7_bid                   ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.bresp   (us7_bresp                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.bvalid  (us7_bvalid                ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.bready  (us7_bready                ), // (axi_master7) => (axi_monitor_m7,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us7_arid                  ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.araddr  (us7_araddr                ), // (axi_master7) => (axi_monitor_m7,bench,bmc300)
	.arlen   (us7_arlen                 ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.arsize  (us7_arsize                ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.arburst (us7_arburst               ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.arlock  ({us7_arlock_b1,us7_arlock}), // () => ()
	.arcache (us7_arcache               ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.arprot  (us7_arprot                ), // (axi_master7) => (axi_monitor_m7,bmc300)
	.arvalid (us7_arvalid               ), // (axi_master7) => (axi_monitor_m7,bench,bmc300)
	.arready (us7_arready               ), // (axi_master7,axi_monitor_m7,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us7_rid                   ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rdata   (us7_rdata                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rresp   (us7_rresp                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rlast   (us7_rlast                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rvalid  (us7_rvalid                ), // (axi_master7,axi_monitor_m7) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us7_rready                )  // (axi_master7) => (axi_monitor_m7,bmc300)
); // end of axi_master7

defparam axi_monitor_m7.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m7.AXI4 = 1'b1;
defparam axi_monitor_m7.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m7.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m7.MASTER_ID = 7;
defparam axi_monitor_m7.SLAVE_ID = 7;
axi_monitor axi_monitor_m7 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us7_awid                  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.awaddr  (us7_awaddr                ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.awlen   (us7_awlen                 ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.awsize  (us7_awsize                ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.awburst (us7_awburst               ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.awlock  ({us7_awlock_b1,us7_awlock}), // () <= ()
	.awcache (us7_awcache               ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.awprot  (us7_awprot                ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.awvalid (us7_awvalid               ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.awready (us7_awready               ), // (axi_master7,axi_monitor_m7,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us7_wid                   ), // (axi_monitor_m7) <= (axi_master7)
	.wdata   (us7_wdata                 ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.wstrb   (us7_wstrb                 ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.wlast   (us7_wlast                 ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.wvalid  (us7_wvalid                ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.wready  (us7_wready                ), // (axi_master7,axi_monitor_m7) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us7_bid                   ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.bresp   (us7_bresp                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.bvalid  (us7_bvalid                ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.bready  (us7_bready                ), // (axi_monitor_m7,bmc300) <= (axi_master7)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us7_arid                  ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.araddr  (us7_araddr                ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.arlen   (us7_arlen                 ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.arsize  (us7_arsize                ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.arburst (us7_arburst               ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.arlock  ({us7_arlock_b1,us7_arlock}), // () <= ()
	.arcache (us7_arcache               ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.arprot  (us7_arprot                ), // (axi_monitor_m7,bmc300) <= (axi_master7)
	.arvalid (us7_arvalid               ), // (axi_monitor_m7,bench,bmc300) <= (axi_master7)
	.arready (us7_arready               ), // (axi_master7,axi_monitor_m7,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us7_rid                   ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rdata   (us7_rdata                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rresp   (us7_rresp                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rlast   (us7_rlast                 ), // (axi_master7,axi_monitor_m7) <= (bmc300)
	.rvalid  (us7_rvalid                ), // (axi_master7,axi_monitor_m7) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us7_rready                )  // (axi_monitor_m7,bmc300) <= (axi_master7)
); // end of axi_monitor_m7

`endif // ATCBMC300_MST7_SUPPORT
`ifdef ATCBMC300_MST8_SUPPORT
defparam axi_master8.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master8.ADDR_START = 0;
defparam axi_master8.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master8.AXI4 = 1'b1;
defparam axi_master8.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master8.DATA_WIDTH = DATA_SIZE;
defparam axi_master8.DELAY_MAX = `ifdef NDS_MST8_DELAY_MAX `NDS_MST8_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master8.ID_WIDTH = US_ID_WIDTH;
defparam axi_master8.MAX_BUF_DEPTH = 256;
defparam axi_master8.MODEL_ID = 8;
defparam axi_master8.TRANS_NUM = `ifdef NDS_MST8_TRANS_NUM `NDS_MST8_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master8.UNALIGN_SUPPORT = 1'b1;
defparam axi_master8.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master8 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us8_awid                  ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.awaddr  (us8_awaddr                ), // (axi_master8) => (axi_monitor_m8,bench,bmc300)
	.awlen   (us8_awlen                 ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.awsize  (us8_awsize                ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.awburst (us8_awburst               ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.awlock  ({us8_awlock_b1,us8_awlock}), // () => ()
	.awcache (us8_awcache               ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.awprot  (us8_awprot                ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.awvalid (us8_awvalid               ), // (axi_master8) => (axi_monitor_m8,bench,bmc300)
	.awready (us8_awready               ), // (axi_master8,axi_monitor_m8,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us8_wid                   ), // (axi_master8) => (axi_monitor_m8)
	.wdata   (us8_wdata                 ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.wstrb   (us8_wstrb                 ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.wlast   (us8_wlast                 ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.wvalid  (us8_wvalid                ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.wready  (us8_wready                ), // (axi_master8,axi_monitor_m8) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us8_bid                   ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.bresp   (us8_bresp                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.bvalid  (us8_bvalid                ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.bready  (us8_bready                ), // (axi_master8) => (axi_monitor_m8,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us8_arid                  ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.araddr  (us8_araddr                ), // (axi_master8) => (axi_monitor_m8,bench,bmc300)
	.arlen   (us8_arlen                 ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.arsize  (us8_arsize                ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.arburst (us8_arburst               ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.arlock  ({us8_arlock_b1,us8_arlock}), // () => ()
	.arcache (us8_arcache               ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.arprot  (us8_arprot                ), // (axi_master8) => (axi_monitor_m8,bmc300)
	.arvalid (us8_arvalid               ), // (axi_master8) => (axi_monitor_m8,bench,bmc300)
	.arready (us8_arready               ), // (axi_master8,axi_monitor_m8,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us8_rid                   ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rdata   (us8_rdata                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rresp   (us8_rresp                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rlast   (us8_rlast                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rvalid  (us8_rvalid                ), // (axi_master8,axi_monitor_m8) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us8_rready                )  // (axi_master8) => (axi_monitor_m8,bmc300)
); // end of axi_master8

defparam axi_monitor_m8.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m8.AXI4 = 1'b1;
defparam axi_monitor_m8.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m8.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m8.MASTER_ID = 8;
defparam axi_monitor_m8.SLAVE_ID = 8;
axi_monitor axi_monitor_m8 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us8_awid                  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.awaddr  (us8_awaddr                ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.awlen   (us8_awlen                 ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.awsize  (us8_awsize                ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.awburst (us8_awburst               ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.awlock  ({us8_awlock_b1,us8_awlock}), // () <= ()
	.awcache (us8_awcache               ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.awprot  (us8_awprot                ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.awvalid (us8_awvalid               ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.awready (us8_awready               ), // (axi_master8,axi_monitor_m8,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us8_wid                   ), // (axi_monitor_m8) <= (axi_master8)
	.wdata   (us8_wdata                 ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.wstrb   (us8_wstrb                 ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.wlast   (us8_wlast                 ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.wvalid  (us8_wvalid                ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.wready  (us8_wready                ), // (axi_master8,axi_monitor_m8) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us8_bid                   ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.bresp   (us8_bresp                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.bvalid  (us8_bvalid                ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.bready  (us8_bready                ), // (axi_monitor_m8,bmc300) <= (axi_master8)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us8_arid                  ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.araddr  (us8_araddr                ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.arlen   (us8_arlen                 ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.arsize  (us8_arsize                ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.arburst (us8_arburst               ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.arlock  ({us8_arlock_b1,us8_arlock}), // () <= ()
	.arcache (us8_arcache               ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.arprot  (us8_arprot                ), // (axi_monitor_m8,bmc300) <= (axi_master8)
	.arvalid (us8_arvalid               ), // (axi_monitor_m8,bench,bmc300) <= (axi_master8)
	.arready (us8_arready               ), // (axi_master8,axi_monitor_m8,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us8_rid                   ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rdata   (us8_rdata                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rresp   (us8_rresp                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rlast   (us8_rlast                 ), // (axi_master8,axi_monitor_m8) <= (bmc300)
	.rvalid  (us8_rvalid                ), // (axi_master8,axi_monitor_m8) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us8_rready                )  // (axi_monitor_m8,bmc300) <= (axi_master8)
); // end of axi_monitor_m8

`endif // ATCBMC300_MST8_SUPPORT
`ifdef ATCBMC300_MST9_SUPPORT
defparam axi_master9.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master9.ADDR_START = 0;
defparam axi_master9.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master9.AXI4 = 1'b1;
defparam axi_master9.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master9.DATA_WIDTH = DATA_SIZE;
defparam axi_master9.DELAY_MAX = `ifdef NDS_MST9_DELAY_MAX `NDS_MST9_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master9.ID_WIDTH = US_ID_WIDTH;
defparam axi_master9.MAX_BUF_DEPTH = 256;
defparam axi_master9.MODEL_ID = 9;
defparam axi_master9.TRANS_NUM = `ifdef NDS_MST9_TRANS_NUM `NDS_MST9_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master9.UNALIGN_SUPPORT = 1'b1;
defparam axi_master9.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master9 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us9_awid                  ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.awaddr  (us9_awaddr                ), // (axi_master9) => (axi_monitor_m9,bench,bmc300)
	.awlen   (us9_awlen                 ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.awsize  (us9_awsize                ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.awburst (us9_awburst               ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.awlock  ({us9_awlock_b1,us9_awlock}), // () => ()
	.awcache (us9_awcache               ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.awprot  (us9_awprot                ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.awvalid (us9_awvalid               ), // (axi_master9) => (axi_monitor_m9,bench,bmc300)
	.awready (us9_awready               ), // (axi_master9,axi_monitor_m9,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us9_wid                   ), // (axi_master9) => (axi_monitor_m9)
	.wdata   (us9_wdata                 ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.wstrb   (us9_wstrb                 ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.wlast   (us9_wlast                 ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.wvalid  (us9_wvalid                ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.wready  (us9_wready                ), // (axi_master9,axi_monitor_m9) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us9_bid                   ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.bresp   (us9_bresp                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.bvalid  (us9_bvalid                ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.bready  (us9_bready                ), // (axi_master9) => (axi_monitor_m9,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us9_arid                  ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.araddr  (us9_araddr                ), // (axi_master9) => (axi_monitor_m9,bench,bmc300)
	.arlen   (us9_arlen                 ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.arsize  (us9_arsize                ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.arburst (us9_arburst               ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.arlock  ({us9_arlock_b1,us9_arlock}), // () => ()
	.arcache (us9_arcache               ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.arprot  (us9_arprot                ), // (axi_master9) => (axi_monitor_m9,bmc300)
	.arvalid (us9_arvalid               ), // (axi_master9) => (axi_monitor_m9,bench,bmc300)
	.arready (us9_arready               ), // (axi_master9,axi_monitor_m9,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us9_rid                   ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rdata   (us9_rdata                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rresp   (us9_rresp                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rlast   (us9_rlast                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rvalid  (us9_rvalid                ), // (axi_master9,axi_monitor_m9) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us9_rready                )  // (axi_master9) => (axi_monitor_m9,bmc300)
); // end of axi_master9

defparam axi_monitor_m9.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m9.AXI4 = 1'b1;
defparam axi_monitor_m9.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m9.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m9.MASTER_ID = 9;
defparam axi_monitor_m9.SLAVE_ID = 9;
axi_monitor axi_monitor_m9 (
	.aclk    (aclk                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                   ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us9_awid                  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.awaddr  (us9_awaddr                ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.awlen   (us9_awlen                 ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.awsize  (us9_awsize                ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.awburst (us9_awburst               ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.awlock  ({us9_awlock_b1,us9_awlock}), // () <= ()
	.awcache (us9_awcache               ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.awprot  (us9_awprot                ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.awvalid (us9_awvalid               ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.awready (us9_awready               ), // (axi_master9,axi_monitor_m9,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us9_wid                   ), // (axi_monitor_m9) <= (axi_master9)
	.wdata   (us9_wdata                 ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.wstrb   (us9_wstrb                 ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.wlast   (us9_wlast                 ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.wvalid  (us9_wvalid                ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.wready  (us9_wready                ), // (axi_master9,axi_monitor_m9) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us9_bid                   ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.bresp   (us9_bresp                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.bvalid  (us9_bvalid                ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.bready  (us9_bready                ), // (axi_monitor_m9,bmc300) <= (axi_master9)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us9_arid                  ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.araddr  (us9_araddr                ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.arlen   (us9_arlen                 ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.arsize  (us9_arsize                ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.arburst (us9_arburst               ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.arlock  ({us9_arlock_b1,us9_arlock}), // () <= ()
	.arcache (us9_arcache               ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.arprot  (us9_arprot                ), // (axi_monitor_m9,bmc300) <= (axi_master9)
	.arvalid (us9_arvalid               ), // (axi_monitor_m9,bench,bmc300) <= (axi_master9)
	.arready (us9_arready               ), // (axi_master9,axi_monitor_m9,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                  ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                     ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us9_rid                   ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rdata   (us9_rdata                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rresp   (us9_rresp                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rlast   (us9_rlast                 ), // (axi_master9,axi_monitor_m9) <= (bmc300)
	.rvalid  (us9_rvalid                ), // (axi_master9,axi_monitor_m9) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us9_rready                )  // (axi_monitor_m9,bmc300) <= (axi_master9)
); // end of axi_monitor_m9

`endif // ATCBMC300_MST9_SUPPORT
`ifdef ATCBMC300_MST10_SUPPORT
defparam axi_master10.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master10.ADDR_START = 0;
defparam axi_master10.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master10.AXI4 = 1'b1;
defparam axi_master10.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master10.DATA_WIDTH = DATA_SIZE;
defparam axi_master10.DELAY_MAX = `ifdef NDS_MST10_DELAY_MAX `NDS_MST10_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master10.ID_WIDTH = US_ID_WIDTH;
defparam axi_master10.MAX_BUF_DEPTH = 256;
defparam axi_master10.MODEL_ID = 10;
defparam axi_master10.TRANS_NUM = `ifdef NDS_MST10_TRANS_NUM `NDS_MST10_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master10.UNALIGN_SUPPORT = 1'b1;
defparam axi_master10.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master10 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us10_awid                   ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.awaddr  (us10_awaddr                 ), // (axi_master10) => (axi_monitor_m10,bench,bmc300)
	.awlen   (us10_awlen                  ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.awsize  (us10_awsize                 ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.awburst (us10_awburst                ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.awlock  ({us10_awlock_b1,us10_awlock}), // () => ()
	.awcache (us10_awcache                ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.awprot  (us10_awprot                 ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.awvalid (us10_awvalid                ), // (axi_master10) => (axi_monitor_m10,bench,bmc300)
	.awready (us10_awready                ), // (axi_master10,axi_monitor_m10,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us10_wid                    ), // (axi_master10) => (axi_monitor_m10)
	.wdata   (us10_wdata                  ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.wstrb   (us10_wstrb                  ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.wlast   (us10_wlast                  ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.wvalid  (us10_wvalid                 ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.wready  (us10_wready                 ), // (axi_master10,axi_monitor_m10) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us10_bid                    ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.bresp   (us10_bresp                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.bvalid  (us10_bvalid                 ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.bready  (us10_bready                 ), // (axi_master10) => (axi_monitor_m10,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us10_arid                   ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.araddr  (us10_araddr                 ), // (axi_master10) => (axi_monitor_m10,bench,bmc300)
	.arlen   (us10_arlen                  ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.arsize  (us10_arsize                 ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.arburst (us10_arburst                ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.arlock  ({us10_arlock_b1,us10_arlock}), // () => ()
	.arcache (us10_arcache                ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.arprot  (us10_arprot                 ), // (axi_master10) => (axi_monitor_m10,bmc300)
	.arvalid (us10_arvalid                ), // (axi_master10) => (axi_monitor_m10,bench,bmc300)
	.arready (us10_arready                ), // (axi_master10,axi_monitor_m10,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us10_rid                    ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rdata   (us10_rdata                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rresp   (us10_rresp                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rlast   (us10_rlast                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rvalid  (us10_rvalid                 ), // (axi_master10,axi_monitor_m10) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us10_rready                 )  // (axi_master10) => (axi_monitor_m10,bmc300)
); // end of axi_master10

defparam axi_monitor_m10.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m10.AXI4 = 1'b1;
defparam axi_monitor_m10.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m10.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m10.MASTER_ID = 10;
defparam axi_monitor_m10.SLAVE_ID = 10;
axi_monitor axi_monitor_m10 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us10_awid                   ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.awaddr  (us10_awaddr                 ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.awlen   (us10_awlen                  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.awsize  (us10_awsize                 ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.awburst (us10_awburst                ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.awlock  ({us10_awlock_b1,us10_awlock}), // () <= ()
	.awcache (us10_awcache                ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.awprot  (us10_awprot                 ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.awvalid (us10_awvalid                ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.awready (us10_awready                ), // (axi_master10,axi_monitor_m10,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us10_wid                    ), // (axi_monitor_m10) <= (axi_master10)
	.wdata   (us10_wdata                  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.wstrb   (us10_wstrb                  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.wlast   (us10_wlast                  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.wvalid  (us10_wvalid                 ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.wready  (us10_wready                 ), // (axi_master10,axi_monitor_m10) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us10_bid                    ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.bresp   (us10_bresp                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.bvalid  (us10_bvalid                 ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.bready  (us10_bready                 ), // (axi_monitor_m10,bmc300) <= (axi_master10)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us10_arid                   ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.araddr  (us10_araddr                 ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.arlen   (us10_arlen                  ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.arsize  (us10_arsize                 ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.arburst (us10_arburst                ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.arlock  ({us10_arlock_b1,us10_arlock}), // () <= ()
	.arcache (us10_arcache                ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.arprot  (us10_arprot                 ), // (axi_monitor_m10,bmc300) <= (axi_master10)
	.arvalid (us10_arvalid                ), // (axi_monitor_m10,bench,bmc300) <= (axi_master10)
	.arready (us10_arready                ), // (axi_master10,axi_monitor_m10,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us10_rid                    ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rdata   (us10_rdata                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rresp   (us10_rresp                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rlast   (us10_rlast                  ), // (axi_master10,axi_monitor_m10) <= (bmc300)
	.rvalid  (us10_rvalid                 ), // (axi_master10,axi_monitor_m10) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us10_rready                 )  // (axi_monitor_m10,bmc300) <= (axi_master10)
); // end of axi_monitor_m10

`endif // ATCBMC300_MST10_SUPPORT
`ifdef ATCBMC300_MST11_SUPPORT
defparam axi_master11.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master11.ADDR_START = 0;
defparam axi_master11.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master11.AXI4 = 1'b1;
defparam axi_master11.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master11.DATA_WIDTH = DATA_SIZE;
defparam axi_master11.DELAY_MAX = `ifdef NDS_MST11_DELAY_MAX `NDS_MST11_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master11.ID_WIDTH = US_ID_WIDTH;
defparam axi_master11.MAX_BUF_DEPTH = 256;
defparam axi_master11.MODEL_ID = 11;
defparam axi_master11.TRANS_NUM = `ifdef NDS_MST11_TRANS_NUM `NDS_MST11_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master11.UNALIGN_SUPPORT = 1'b1;
defparam axi_master11.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master11 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us11_awid                   ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.awaddr  (us11_awaddr                 ), // (axi_master11) => (axi_monitor_m11,bench,bmc300)
	.awlen   (us11_awlen                  ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.awsize  (us11_awsize                 ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.awburst (us11_awburst                ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.awlock  ({us11_awlock_b1,us11_awlock}), // () => ()
	.awcache (us11_awcache                ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.awprot  (us11_awprot                 ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.awvalid (us11_awvalid                ), // (axi_master11) => (axi_monitor_m11,bench,bmc300)
	.awready (us11_awready                ), // (axi_master11,axi_monitor_m11,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us11_wid                    ), // (axi_master11) => (axi_monitor_m11)
	.wdata   (us11_wdata                  ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.wstrb   (us11_wstrb                  ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.wlast   (us11_wlast                  ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.wvalid  (us11_wvalid                 ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.wready  (us11_wready                 ), // (axi_master11,axi_monitor_m11) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us11_bid                    ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.bresp   (us11_bresp                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.bvalid  (us11_bvalid                 ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.bready  (us11_bready                 ), // (axi_master11) => (axi_monitor_m11,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us11_arid                   ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.araddr  (us11_araddr                 ), // (axi_master11) => (axi_monitor_m11,bench,bmc300)
	.arlen   (us11_arlen                  ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.arsize  (us11_arsize                 ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.arburst (us11_arburst                ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.arlock  ({us11_arlock_b1,us11_arlock}), // () => ()
	.arcache (us11_arcache                ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.arprot  (us11_arprot                 ), // (axi_master11) => (axi_monitor_m11,bmc300)
	.arvalid (us11_arvalid                ), // (axi_master11) => (axi_monitor_m11,bench,bmc300)
	.arready (us11_arready                ), // (axi_master11,axi_monitor_m11,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us11_rid                    ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rdata   (us11_rdata                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rresp   (us11_rresp                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rlast   (us11_rlast                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rvalid  (us11_rvalid                 ), // (axi_master11,axi_monitor_m11) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us11_rready                 )  // (axi_master11) => (axi_monitor_m11,bmc300)
); // end of axi_master11

defparam axi_monitor_m11.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m11.AXI4 = 1'b1;
defparam axi_monitor_m11.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m11.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m11.MASTER_ID = 11;
defparam axi_monitor_m11.SLAVE_ID = 11;
axi_monitor axi_monitor_m11 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us11_awid                   ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.awaddr  (us11_awaddr                 ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.awlen   (us11_awlen                  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.awsize  (us11_awsize                 ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.awburst (us11_awburst                ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.awlock  ({us11_awlock_b1,us11_awlock}), // () <= ()
	.awcache (us11_awcache                ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.awprot  (us11_awprot                 ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.awvalid (us11_awvalid                ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.awready (us11_awready                ), // (axi_master11,axi_monitor_m11,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us11_wid                    ), // (axi_monitor_m11) <= (axi_master11)
	.wdata   (us11_wdata                  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.wstrb   (us11_wstrb                  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.wlast   (us11_wlast                  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.wvalid  (us11_wvalid                 ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.wready  (us11_wready                 ), // (axi_master11,axi_monitor_m11) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us11_bid                    ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.bresp   (us11_bresp                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.bvalid  (us11_bvalid                 ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.bready  (us11_bready                 ), // (axi_monitor_m11,bmc300) <= (axi_master11)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us11_arid                   ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.araddr  (us11_araddr                 ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.arlen   (us11_arlen                  ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.arsize  (us11_arsize                 ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.arburst (us11_arburst                ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.arlock  ({us11_arlock_b1,us11_arlock}), // () <= ()
	.arcache (us11_arcache                ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.arprot  (us11_arprot                 ), // (axi_monitor_m11,bmc300) <= (axi_master11)
	.arvalid (us11_arvalid                ), // (axi_monitor_m11,bench,bmc300) <= (axi_master11)
	.arready (us11_arready                ), // (axi_master11,axi_monitor_m11,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us11_rid                    ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rdata   (us11_rdata                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rresp   (us11_rresp                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rlast   (us11_rlast                  ), // (axi_master11,axi_monitor_m11) <= (bmc300)
	.rvalid  (us11_rvalid                 ), // (axi_master11,axi_monitor_m11) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us11_rready                 )  // (axi_monitor_m11,bmc300) <= (axi_master11)
); // end of axi_monitor_m11

`endif // ATCBMC300_MST11_SUPPORT
`ifdef ATCBMC300_MST12_SUPPORT
defparam axi_master12.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master12.ADDR_START = 0;
defparam axi_master12.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master12.AXI4 = 1'b1;
defparam axi_master12.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master12.DATA_WIDTH = DATA_SIZE;
defparam axi_master12.DELAY_MAX = `ifdef NDS_MST12_DELAY_MAX `NDS_MST12_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master12.ID_WIDTH = US_ID_WIDTH;
defparam axi_master12.MAX_BUF_DEPTH = 256;
defparam axi_master12.MODEL_ID = 12;
defparam axi_master12.TRANS_NUM = `ifdef NDS_MST12_TRANS_NUM `NDS_MST12_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master12.UNALIGN_SUPPORT = 1'b1;
defparam axi_master12.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master12 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us12_awid                   ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.awaddr  (us12_awaddr                 ), // (axi_master12) => (axi_monitor_m12,bench,bmc300)
	.awlen   (us12_awlen                  ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.awsize  (us12_awsize                 ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.awburst (us12_awburst                ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.awlock  ({us12_awlock_b1,us12_awlock}), // () => ()
	.awcache (us12_awcache                ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.awprot  (us12_awprot                 ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.awvalid (us12_awvalid                ), // (axi_master12) => (axi_monitor_m12,bench,bmc300)
	.awready (us12_awready                ), // (axi_master12,axi_monitor_m12,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us12_wid                    ), // (axi_master12) => (axi_monitor_m12)
	.wdata   (us12_wdata                  ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.wstrb   (us12_wstrb                  ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.wlast   (us12_wlast                  ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.wvalid  (us12_wvalid                 ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.wready  (us12_wready                 ), // (axi_master12,axi_monitor_m12) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us12_bid                    ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.bresp   (us12_bresp                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.bvalid  (us12_bvalid                 ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.bready  (us12_bready                 ), // (axi_master12) => (axi_monitor_m12,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us12_arid                   ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.araddr  (us12_araddr                 ), // (axi_master12) => (axi_monitor_m12,bench,bmc300)
	.arlen   (us12_arlen                  ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.arsize  (us12_arsize                 ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.arburst (us12_arburst                ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.arlock  ({us12_arlock_b1,us12_arlock}), // () => ()
	.arcache (us12_arcache                ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.arprot  (us12_arprot                 ), // (axi_master12) => (axi_monitor_m12,bmc300)
	.arvalid (us12_arvalid                ), // (axi_master12) => (axi_monitor_m12,bench,bmc300)
	.arready (us12_arready                ), // (axi_master12,axi_monitor_m12,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us12_rid                    ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rdata   (us12_rdata                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rresp   (us12_rresp                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rlast   (us12_rlast                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rvalid  (us12_rvalid                 ), // (axi_master12,axi_monitor_m12) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us12_rready                 )  // (axi_master12) => (axi_monitor_m12,bmc300)
); // end of axi_master12

defparam axi_monitor_m12.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m12.AXI4 = 1'b1;
defparam axi_monitor_m12.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m12.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m12.MASTER_ID = 12;
defparam axi_monitor_m12.SLAVE_ID = 12;
axi_monitor axi_monitor_m12 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us12_awid                   ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.awaddr  (us12_awaddr                 ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.awlen   (us12_awlen                  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.awsize  (us12_awsize                 ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.awburst (us12_awburst                ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.awlock  ({us12_awlock_b1,us12_awlock}), // () <= ()
	.awcache (us12_awcache                ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.awprot  (us12_awprot                 ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.awvalid (us12_awvalid                ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.awready (us12_awready                ), // (axi_master12,axi_monitor_m12,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us12_wid                    ), // (axi_monitor_m12) <= (axi_master12)
	.wdata   (us12_wdata                  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.wstrb   (us12_wstrb                  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.wlast   (us12_wlast                  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.wvalid  (us12_wvalid                 ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.wready  (us12_wready                 ), // (axi_master12,axi_monitor_m12) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us12_bid                    ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.bresp   (us12_bresp                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.bvalid  (us12_bvalid                 ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.bready  (us12_bready                 ), // (axi_monitor_m12,bmc300) <= (axi_master12)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us12_arid                   ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.araddr  (us12_araddr                 ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.arlen   (us12_arlen                  ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.arsize  (us12_arsize                 ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.arburst (us12_arburst                ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.arlock  ({us12_arlock_b1,us12_arlock}), // () <= ()
	.arcache (us12_arcache                ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.arprot  (us12_arprot                 ), // (axi_monitor_m12,bmc300) <= (axi_master12)
	.arvalid (us12_arvalid                ), // (axi_monitor_m12,bench,bmc300) <= (axi_master12)
	.arready (us12_arready                ), // (axi_master12,axi_monitor_m12,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us12_rid                    ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rdata   (us12_rdata                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rresp   (us12_rresp                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rlast   (us12_rlast                  ), // (axi_master12,axi_monitor_m12) <= (bmc300)
	.rvalid  (us12_rvalid                 ), // (axi_master12,axi_monitor_m12) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us12_rready                 )  // (axi_monitor_m12,bmc300) <= (axi_master12)
); // end of axi_monitor_m12

`endif // ATCBMC300_MST12_SUPPORT
`ifdef ATCBMC300_MST13_SUPPORT
defparam axi_master13.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master13.ADDR_START = 0;
defparam axi_master13.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master13.AXI4 = 1'b1;
defparam axi_master13.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master13.DATA_WIDTH = DATA_SIZE;
defparam axi_master13.DELAY_MAX = `ifdef NDS_MST13_DELAY_MAX `NDS_MST13_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master13.ID_WIDTH = US_ID_WIDTH;
defparam axi_master13.MAX_BUF_DEPTH = 256;
defparam axi_master13.MODEL_ID = 13;
defparam axi_master13.TRANS_NUM = `ifdef NDS_MST13_TRANS_NUM `NDS_MST13_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master13.UNALIGN_SUPPORT = 1'b1;
defparam axi_master13.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master13 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us13_awid                   ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.awaddr  (us13_awaddr                 ), // (axi_master13) => (axi_monitor_m13,bench,bmc300)
	.awlen   (us13_awlen                  ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.awsize  (us13_awsize                 ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.awburst (us13_awburst                ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.awlock  ({us13_awlock_b1,us13_awlock}), // () => ()
	.awcache (us13_awcache                ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.awprot  (us13_awprot                 ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.awvalid (us13_awvalid                ), // (axi_master13) => (axi_monitor_m13,bench,bmc300)
	.awready (us13_awready                ), // (axi_master13,axi_monitor_m13,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us13_wid                    ), // (axi_master13) => (axi_monitor_m13)
	.wdata   (us13_wdata                  ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.wstrb   (us13_wstrb                  ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.wlast   (us13_wlast                  ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.wvalid  (us13_wvalid                 ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.wready  (us13_wready                 ), // (axi_master13,axi_monitor_m13) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us13_bid                    ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.bresp   (us13_bresp                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.bvalid  (us13_bvalid                 ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.bready  (us13_bready                 ), // (axi_master13) => (axi_monitor_m13,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us13_arid                   ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.araddr  (us13_araddr                 ), // (axi_master13) => (axi_monitor_m13,bench,bmc300)
	.arlen   (us13_arlen                  ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.arsize  (us13_arsize                 ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.arburst (us13_arburst                ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.arlock  ({us13_arlock_b1,us13_arlock}), // () => ()
	.arcache (us13_arcache                ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.arprot  (us13_arprot                 ), // (axi_master13) => (axi_monitor_m13,bmc300)
	.arvalid (us13_arvalid                ), // (axi_master13) => (axi_monitor_m13,bench,bmc300)
	.arready (us13_arready                ), // (axi_master13,axi_monitor_m13,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us13_rid                    ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rdata   (us13_rdata                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rresp   (us13_rresp                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rlast   (us13_rlast                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rvalid  (us13_rvalid                 ), // (axi_master13,axi_monitor_m13) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us13_rready                 )  // (axi_master13) => (axi_monitor_m13,bmc300)
); // end of axi_master13

defparam axi_monitor_m13.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m13.AXI4 = 1'b1;
defparam axi_monitor_m13.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m13.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m13.MASTER_ID = 13;
defparam axi_monitor_m13.SLAVE_ID = 13;
axi_monitor axi_monitor_m13 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us13_awid                   ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.awaddr  (us13_awaddr                 ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.awlen   (us13_awlen                  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.awsize  (us13_awsize                 ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.awburst (us13_awburst                ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.awlock  ({us13_awlock_b1,us13_awlock}), // () <= ()
	.awcache (us13_awcache                ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.awprot  (us13_awprot                 ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.awvalid (us13_awvalid                ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.awready (us13_awready                ), // (axi_master13,axi_monitor_m13,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us13_wid                    ), // (axi_monitor_m13) <= (axi_master13)
	.wdata   (us13_wdata                  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.wstrb   (us13_wstrb                  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.wlast   (us13_wlast                  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.wvalid  (us13_wvalid                 ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.wready  (us13_wready                 ), // (axi_master13,axi_monitor_m13) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us13_bid                    ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.bresp   (us13_bresp                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.bvalid  (us13_bvalid                 ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.bready  (us13_bready                 ), // (axi_monitor_m13,bmc300) <= (axi_master13)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us13_arid                   ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.araddr  (us13_araddr                 ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.arlen   (us13_arlen                  ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.arsize  (us13_arsize                 ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.arburst (us13_arburst                ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.arlock  ({us13_arlock_b1,us13_arlock}), // () <= ()
	.arcache (us13_arcache                ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.arprot  (us13_arprot                 ), // (axi_monitor_m13,bmc300) <= (axi_master13)
	.arvalid (us13_arvalid                ), // (axi_monitor_m13,bench,bmc300) <= (axi_master13)
	.arready (us13_arready                ), // (axi_master13,axi_monitor_m13,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us13_rid                    ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rdata   (us13_rdata                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rresp   (us13_rresp                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rlast   (us13_rlast                  ), // (axi_master13,axi_monitor_m13) <= (bmc300)
	.rvalid  (us13_rvalid                 ), // (axi_master13,axi_monitor_m13) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us13_rready                 )  // (axi_monitor_m13,bmc300) <= (axi_master13)
); // end of axi_monitor_m13

`endif // ATCBMC300_MST13_SUPPORT
`ifdef ATCBMC300_MST14_SUPPORT
defparam axi_master14.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master14.ADDR_START = 0;
defparam axi_master14.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master14.AXI4 = 1'b1;
defparam axi_master14.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master14.DATA_WIDTH = DATA_SIZE;
defparam axi_master14.DELAY_MAX = `ifdef NDS_MST14_DELAY_MAX `NDS_MST14_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master14.ID_WIDTH = US_ID_WIDTH;
defparam axi_master14.MAX_BUF_DEPTH = 256;
defparam axi_master14.MODEL_ID = 14;
defparam axi_master14.TRANS_NUM = `ifdef NDS_MST14_TRANS_NUM `NDS_MST14_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master14.UNALIGN_SUPPORT = 1'b1;
defparam axi_master14.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master14 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us14_awid                   ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.awaddr  (us14_awaddr                 ), // (axi_master14) => (axi_monitor_m14,bench,bmc300)
	.awlen   (us14_awlen                  ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.awsize  (us14_awsize                 ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.awburst (us14_awburst                ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.awlock  ({us14_awlock_b1,us14_awlock}), // () => ()
	.awcache (us14_awcache                ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.awprot  (us14_awprot                 ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.awvalid (us14_awvalid                ), // (axi_master14) => (axi_monitor_m14,bench,bmc300)
	.awready (us14_awready                ), // (axi_master14,axi_monitor_m14,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us14_wid                    ), // (axi_master14) => (axi_monitor_m14)
	.wdata   (us14_wdata                  ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.wstrb   (us14_wstrb                  ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.wlast   (us14_wlast                  ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.wvalid  (us14_wvalid                 ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.wready  (us14_wready                 ), // (axi_master14,axi_monitor_m14) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us14_bid                    ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.bresp   (us14_bresp                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.bvalid  (us14_bvalid                 ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.bready  (us14_bready                 ), // (axi_master14) => (axi_monitor_m14,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us14_arid                   ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.araddr  (us14_araddr                 ), // (axi_master14) => (axi_monitor_m14,bench,bmc300)
	.arlen   (us14_arlen                  ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.arsize  (us14_arsize                 ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.arburst (us14_arburst                ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.arlock  ({us14_arlock_b1,us14_arlock}), // () => ()
	.arcache (us14_arcache                ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.arprot  (us14_arprot                 ), // (axi_master14) => (axi_monitor_m14,bmc300)
	.arvalid (us14_arvalid                ), // (axi_master14) => (axi_monitor_m14,bench,bmc300)
	.arready (us14_arready                ), // (axi_master14,axi_monitor_m14,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us14_rid                    ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rdata   (us14_rdata                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rresp   (us14_rresp                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rlast   (us14_rlast                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rvalid  (us14_rvalid                 ), // (axi_master14,axi_monitor_m14) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us14_rready                 )  // (axi_master14) => (axi_monitor_m14,bmc300)
); // end of axi_master14

defparam axi_monitor_m14.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m14.AXI4 = 1'b1;
defparam axi_monitor_m14.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m14.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m14.MASTER_ID = 14;
defparam axi_monitor_m14.SLAVE_ID = 14;
axi_monitor axi_monitor_m14 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us14_awid                   ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.awaddr  (us14_awaddr                 ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.awlen   (us14_awlen                  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.awsize  (us14_awsize                 ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.awburst (us14_awburst                ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.awlock  ({us14_awlock_b1,us14_awlock}), // () <= ()
	.awcache (us14_awcache                ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.awprot  (us14_awprot                 ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.awvalid (us14_awvalid                ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.awready (us14_awready                ), // (axi_master14,axi_monitor_m14,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us14_wid                    ), // (axi_monitor_m14) <= (axi_master14)
	.wdata   (us14_wdata                  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.wstrb   (us14_wstrb                  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.wlast   (us14_wlast                  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.wvalid  (us14_wvalid                 ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.wready  (us14_wready                 ), // (axi_master14,axi_monitor_m14) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us14_bid                    ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.bresp   (us14_bresp                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.bvalid  (us14_bvalid                 ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.bready  (us14_bready                 ), // (axi_monitor_m14,bmc300) <= (axi_master14)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us14_arid                   ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.araddr  (us14_araddr                 ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.arlen   (us14_arlen                  ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.arsize  (us14_arsize                 ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.arburst (us14_arburst                ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.arlock  ({us14_arlock_b1,us14_arlock}), // () <= ()
	.arcache (us14_arcache                ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.arprot  (us14_arprot                 ), // (axi_monitor_m14,bmc300) <= (axi_master14)
	.arvalid (us14_arvalid                ), // (axi_monitor_m14,bench,bmc300) <= (axi_master14)
	.arready (us14_arready                ), // (axi_master14,axi_monitor_m14,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us14_rid                    ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rdata   (us14_rdata                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rresp   (us14_rresp                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rlast   (us14_rlast                  ), // (axi_master14,axi_monitor_m14) <= (bmc300)
	.rvalid  (us14_rvalid                 ), // (axi_master14,axi_monitor_m14) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us14_rready                 )  // (axi_monitor_m14,bmc300) <= (axi_master14)
); // end of axi_monitor_m14

`endif // ATCBMC300_MST14_SUPPORT
`ifdef ATCBMC300_MST15_SUPPORT
defparam axi_master15.ADDR_SIZE = (1<<ADDR_WIDTH);
defparam axi_master15.ADDR_START = 0;
defparam axi_master15.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_master15.AXI4 = 1'b1;
defparam axi_master15.AXI4_AXLEN_LT16 = 1'b0;
defparam axi_master15.DATA_WIDTH = DATA_SIZE;
defparam axi_master15.DELAY_MAX = `ifdef NDS_MST15_DELAY_MAX `NDS_MST15_DELAY_MAX `else `NDS_DEFAULT_DELAY_MAX `endif;
defparam axi_master15.ID_WIDTH = US_ID_WIDTH;
defparam axi_master15.MAX_BUF_DEPTH = 256;
defparam axi_master15.MODEL_ID = 15;
defparam axi_master15.TRANS_NUM = `ifdef NDS_MST15_TRANS_NUM `NDS_MST15_TRANS_NUM `else `NDS_DEFAULT_TRANS_NUM `endif;
defparam axi_master15.UNALIGN_SUPPORT = 1'b1;
defparam axi_master15.WAIT_TIMEOUT_CNT = 1000000;
axi_master_model axi_master15 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us15_awid                   ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.awaddr  (us15_awaddr                 ), // (axi_master15) => (axi_monitor_m15,bench,bmc300)
	.awlen   (us15_awlen                  ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.awsize  (us15_awsize                 ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.awburst (us15_awburst                ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.awlock  ({us15_awlock_b1,us15_awlock}), // () => ()
	.awcache (us15_awcache                ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.awprot  (us15_awprot                 ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.awvalid (us15_awvalid                ), // (axi_master15) => (axi_monitor_m15,bench,bmc300)
	.awready (us15_awready                ), // (axi_master15,axi_monitor_m15,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us15_wid                    ), // (axi_master15) => (axi_monitor_m15)
	.wdata   (us15_wdata                  ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.wstrb   (us15_wstrb                  ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.wlast   (us15_wlast                  ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.wvalid  (us15_wvalid                 ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.wready  (us15_wready                 ), // (axi_master15,axi_monitor_m15) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us15_bid                    ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.bresp   (us15_bresp                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.bvalid  (us15_bvalid                 ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.bready  (us15_bready                 ), // (axi_master15) => (axi_monitor_m15,bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us15_arid                   ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.araddr  (us15_araddr                 ), // (axi_master15) => (axi_monitor_m15,bench,bmc300)
	.arlen   (us15_arlen                  ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.arsize  (us15_arsize                 ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.arburst (us15_arburst                ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.arlock  ({us15_arlock_b1,us15_arlock}), // () => ()
	.arcache (us15_arcache                ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.arprot  (us15_arprot                 ), // (axi_master15) => (axi_monitor_m15,bmc300)
	.arvalid (us15_arvalid                ), // (axi_master15) => (axi_monitor_m15,bench,bmc300)
	.arready (us15_arready                ), // (axi_master15,axi_monitor_m15,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9) => (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us15_rid                    ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rdata   (us15_rdata                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rresp   (us15_rresp                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rlast   (us15_rlast                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rvalid  (us15_rvalid                 ), // (axi_master15,axi_monitor_m15) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us15_rready                 )  // (axi_master15) => (axi_monitor_m15,bmc300)
); // end of axi_master15

defparam axi_monitor_m15.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_m15.AXI4 = 1'b1;
defparam axi_monitor_m15.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_m15.ID_WIDTH = US_ID_WIDTH;
defparam axi_monitor_m15.MASTER_ID = 15;
defparam axi_monitor_m15.SLAVE_ID = 15;
axi_monitor axi_monitor_m15 (
	.aclk    (aclk                        ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn                     ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (us15_awid                   ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.awaddr  (us15_awaddr                 ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.awlen   (us15_awlen                  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.awsize  (us15_awsize                 ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.awburst (us15_awburst                ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.awlock  ({us15_awlock_b1,us15_awlock}), // () <= ()
	.awcache (us15_awcache                ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.awprot  (us15_awprot                 ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.awvalid (us15_awvalid                ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.awready (us15_awready                ), // (axi_master15,axi_monitor_m15,bench) <= (bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (us15_wid                    ), // (axi_monitor_m15) <= (axi_master15)
	.wdata   (us15_wdata                  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.wstrb   (us15_wstrb                  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.wlast   (us15_wlast                  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.wvalid  (us15_wvalid                 ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.wready  (us15_wready                 ), // (axi_master15,axi_monitor_m15) <= (bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (us15_bid                    ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.bresp   (us15_bresp                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.bvalid  (us15_bvalid                 ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.bready  (us15_bready                 ), // (axi_monitor_m15,bmc300) <= (axi_master15)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (us15_arid                   ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.araddr  (us15_araddr                 ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.arlen   (us15_arlen                  ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.arsize  (us15_arsize                 ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.arburst (us15_arburst                ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.arlock  ({us15_arlock_b1,us15_arlock}), // () <= ()
	.arcache (us15_arcache                ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.arprot  (us15_arprot                 ), // (axi_monitor_m15,bmc300) <= (axi_master15)
	.arvalid (us15_arvalid                ), // (axi_monitor_m15,bench,bmc300) <= (axi_master15)
	.arready (us15_arready                ), // (axi_master15,axi_monitor_m15,bench) <= (bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion                    ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos                       ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser                      ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (us15_rid                    ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rdata   (us15_rdata                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rresp   (us15_rresp                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rlast   (us15_rlast                  ), // (axi_master15,axi_monitor_m15) <= (bmc300)
	.rvalid  (us15_rvalid                 ), // (axi_master15,axi_monitor_m15) <= (bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser                       ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (us15_rready                 )  // (axi_monitor_m15,bmc300) <= (axi_master15)
); // end of axi_monitor_m15

`endif // ATCBMC300_MST15_SUPPORT
`ifdef ATCBMC300_SLV1_SUPPORT
defparam axi_slave1.ADDR_DECODE_WIDTH = `ATCBMC300_SLV1_SIZE+19;
defparam axi_slave1.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave1.AXI4 = 1'b1;
defparam axi_slave1.DATA_WIDTH = DATA_SIZE;
defparam axi_slave1.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave1.MEM_ADDR_WIDTH = `ATCBMC300_SLV1_SIZE+19;
defparam axi_slave1.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave1 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds1_awid         ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awaddr  (ds1_awaddr       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awlen   (ds1_awlen        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awsize  (ds1_awsize       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awburst (ds1_awburst      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awlock  ({1'b0,ds1_awlock}), // () <= ()
	.awcache (ds1_awcache      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awprot  (ds1_awprot       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awvalid (ds1_awvalid      ), // (axi_monitor_s1,axi_slave1,bench) <= (bmc300)
	.awready (ds1_awready      ), // (axi_slave1) => (axi_monitor_s1,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds1_wid          ), // (axi_monitor_s1,axi_slave1) <= ()
	.wdata   (ds1_wdata        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wstrb   (ds1_wstrb        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wlast   (ds1_wlast        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wvalid  (ds1_wvalid       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wready  (ds1_wready       ), // (axi_slave1) => (axi_monitor_s1,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds1_bid          ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.bresp   (ds1_bresp        ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.bvalid  (ds1_bvalid       ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.bready  (ds1_bready       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds1_arid         ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.araddr  (ds1_araddr       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arlen   (ds1_arlen        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arsize  (ds1_arsize       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arburst (ds1_arburst      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arlock  ({1'b0,ds1_arlock}), // () <= ()
	.arcache (ds1_arcache      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arprot  (ds1_arprot       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arvalid (ds1_arvalid      ), // (axi_monitor_s1,axi_slave1,bench) <= (bmc300)
	.arready (ds1_arready      ), // (axi_slave1) => (axi_monitor_s1,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds1_rid          ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.rdata   (ds1_rdata        ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.rresp   (ds1_rresp        ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.rlast   (ds1_rlast        ), // (axi_slave1) => (axi_monitor_s1,bmc300)
	.rvalid  (ds1_rvalid       ), // (axi_slave1) => (axi_monitor_s1,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds1_rready       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave1) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave1

defparam axi_monitor_s1.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s1.AXI4 = 1'b1;
defparam axi_monitor_s1.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s1.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s1.MASTER_ID = 101;
defparam axi_monitor_s1.SLAVE_ID = 101;
axi_monitor axi_monitor_s1 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds1_awid         ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awaddr  (ds1_awaddr       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awlen   (ds1_awlen        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awsize  (ds1_awsize       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awburst (ds1_awburst      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awlock  ({1'b0,ds1_awlock}), // () <= ()
	.awcache (ds1_awcache      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awprot  (ds1_awprot       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.awvalid (ds1_awvalid      ), // (axi_monitor_s1,axi_slave1,bench) <= (bmc300)
	.awready (ds1_awready      ), // (axi_monitor_s1,bench,bmc300) <= (axi_slave1)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds1_wid          ), // (axi_monitor_s1,axi_slave1) <= ()
	.wdata   (ds1_wdata        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wstrb   (ds1_wstrb        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wlast   (ds1_wlast        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wvalid  (ds1_wvalid       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.wready  (ds1_wready       ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds1_bid          ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.bresp   (ds1_bresp        ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.bvalid  (ds1_bvalid       ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.bready  (ds1_bready       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds1_arid         ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.araddr  (ds1_araddr       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arlen   (ds1_arlen        ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arsize  (ds1_arsize       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arburst (ds1_arburst      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arlock  ({1'b0,ds1_arlock}), // () <= ()
	.arcache (ds1_arcache      ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arprot  (ds1_arprot       ), // (axi_monitor_s1,axi_slave1) <= (bmc300)
	.arvalid (ds1_arvalid      ), // (axi_monitor_s1,axi_slave1,bench) <= (bmc300)
	.arready (ds1_arready      ), // (axi_monitor_s1,bench,bmc300) <= (axi_slave1)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds1_rid          ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.rdata   (ds1_rdata        ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.rresp   (ds1_rresp        ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.rlast   (ds1_rlast        ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
	.rvalid  (ds1_rvalid       ), // (axi_monitor_s1,bmc300) <= (axi_slave1)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds1_rready       )  // (axi_monitor_s1,axi_slave1) <= (bmc300)
); // end of axi_monitor_s1

`endif // ATCBMC300_SLV1_SUPPORT
`ifdef ATCBMC300_SLV2_SUPPORT
defparam axi_slave2.ADDR_DECODE_WIDTH = `ATCBMC300_SLV2_SIZE+19;
defparam axi_slave2.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave2.AXI4 = 1'b1;
defparam axi_slave2.DATA_WIDTH = DATA_SIZE;
defparam axi_slave2.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave2.MEM_ADDR_WIDTH = `ATCBMC300_SLV2_SIZE+19;
defparam axi_slave2.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave2 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds2_awid         ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awaddr  (ds2_awaddr       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awlen   (ds2_awlen        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awsize  (ds2_awsize       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awburst (ds2_awburst      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awlock  ({1'b0,ds2_awlock}), // () <= ()
	.awcache (ds2_awcache      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awprot  (ds2_awprot       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awvalid (ds2_awvalid      ), // (axi_monitor_s2,axi_slave2,bench) <= (bmc300)
	.awready (ds2_awready      ), // (axi_slave2) => (axi_monitor_s2,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds2_wid          ), // (axi_monitor_s2,axi_slave2) <= ()
	.wdata   (ds2_wdata        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wstrb   (ds2_wstrb        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wlast   (ds2_wlast        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wvalid  (ds2_wvalid       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wready  (ds2_wready       ), // (axi_slave2) => (axi_monitor_s2,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds2_bid          ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.bresp   (ds2_bresp        ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.bvalid  (ds2_bvalid       ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.bready  (ds2_bready       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds2_arid         ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.araddr  (ds2_araddr       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arlen   (ds2_arlen        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arsize  (ds2_arsize       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arburst (ds2_arburst      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arlock  ({1'b0,ds2_arlock}), // () <= ()
	.arcache (ds2_arcache      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arprot  (ds2_arprot       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arvalid (ds2_arvalid      ), // (axi_monitor_s2,axi_slave2,bench) <= (bmc300)
	.arready (ds2_arready      ), // (axi_slave2) => (axi_monitor_s2,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds2_rid          ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.rdata   (ds2_rdata        ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.rresp   (ds2_rresp        ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.rlast   (ds2_rlast        ), // (axi_slave2) => (axi_monitor_s2,bmc300)
	.rvalid  (ds2_rvalid       ), // (axi_slave2) => (axi_monitor_s2,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds2_rready       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave2) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave2

defparam axi_monitor_s2.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s2.AXI4 = 1'b1;
defparam axi_monitor_s2.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s2.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s2.MASTER_ID = 102;
defparam axi_monitor_s2.SLAVE_ID = 102;
axi_monitor axi_monitor_s2 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds2_awid         ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awaddr  (ds2_awaddr       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awlen   (ds2_awlen        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awsize  (ds2_awsize       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awburst (ds2_awburst      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awlock  ({1'b0,ds2_awlock}), // () <= ()
	.awcache (ds2_awcache      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awprot  (ds2_awprot       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.awvalid (ds2_awvalid      ), // (axi_monitor_s2,axi_slave2,bench) <= (bmc300)
	.awready (ds2_awready      ), // (axi_monitor_s2,bench,bmc300) <= (axi_slave2)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds2_wid          ), // (axi_monitor_s2,axi_slave2) <= ()
	.wdata   (ds2_wdata        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wstrb   (ds2_wstrb        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wlast   (ds2_wlast        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wvalid  (ds2_wvalid       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.wready  (ds2_wready       ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds2_bid          ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.bresp   (ds2_bresp        ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.bvalid  (ds2_bvalid       ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.bready  (ds2_bready       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds2_arid         ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.araddr  (ds2_araddr       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arlen   (ds2_arlen        ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arsize  (ds2_arsize       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arburst (ds2_arburst      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arlock  ({1'b0,ds2_arlock}), // () <= ()
	.arcache (ds2_arcache      ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arprot  (ds2_arprot       ), // (axi_monitor_s2,axi_slave2) <= (bmc300)
	.arvalid (ds2_arvalid      ), // (axi_monitor_s2,axi_slave2,bench) <= (bmc300)
	.arready (ds2_arready      ), // (axi_monitor_s2,bench,bmc300) <= (axi_slave2)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds2_rid          ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.rdata   (ds2_rdata        ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.rresp   (ds2_rresp        ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.rlast   (ds2_rlast        ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
	.rvalid  (ds2_rvalid       ), // (axi_monitor_s2,bmc300) <= (axi_slave2)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds2_rready       )  // (axi_monitor_s2,axi_slave2) <= (bmc300)
); // end of axi_monitor_s2

`endif // ATCBMC300_SLV2_SUPPORT
`ifdef ATCBMC300_SLV3_SUPPORT
defparam axi_slave3.ADDR_DECODE_WIDTH = `ATCBMC300_SLV3_SIZE+19;
defparam axi_slave3.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave3.AXI4 = 1'b1;
defparam axi_slave3.DATA_WIDTH = DATA_SIZE;
defparam axi_slave3.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave3.MEM_ADDR_WIDTH = `ATCBMC300_SLV3_SIZE+19;
defparam axi_slave3.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave3 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds3_awid         ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awaddr  (ds3_awaddr       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awlen   (ds3_awlen        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awsize  (ds3_awsize       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awburst (ds3_awburst      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awlock  ({1'b0,ds3_awlock}), // () <= ()
	.awcache (ds3_awcache      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awprot  (ds3_awprot       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awvalid (ds3_awvalid      ), // (axi_monitor_s3,axi_slave3,bench) <= (bmc300)
	.awready (ds3_awready      ), // (axi_slave3) => (axi_monitor_s3,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds3_wid          ), // (axi_monitor_s3,axi_slave3) <= ()
	.wdata   (ds3_wdata        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wstrb   (ds3_wstrb        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wlast   (ds3_wlast        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wvalid  (ds3_wvalid       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wready  (ds3_wready       ), // (axi_slave3) => (axi_monitor_s3,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds3_bid          ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.bresp   (ds3_bresp        ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.bvalid  (ds3_bvalid       ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.bready  (ds3_bready       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds3_arid         ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.araddr  (ds3_araddr       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arlen   (ds3_arlen        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arsize  (ds3_arsize       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arburst (ds3_arburst      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arlock  ({1'b0,ds3_arlock}), // () <= ()
	.arcache (ds3_arcache      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arprot  (ds3_arprot       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arvalid (ds3_arvalid      ), // (axi_monitor_s3,axi_slave3,bench) <= (bmc300)
	.arready (ds3_arready      ), // (axi_slave3) => (axi_monitor_s3,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds3_rid          ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.rdata   (ds3_rdata        ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.rresp   (ds3_rresp        ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.rlast   (ds3_rlast        ), // (axi_slave3) => (axi_monitor_s3,bmc300)
	.rvalid  (ds3_rvalid       ), // (axi_slave3) => (axi_monitor_s3,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds3_rready       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave3) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave3

defparam axi_monitor_s3.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s3.AXI4 = 1'b1;
defparam axi_monitor_s3.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s3.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s3.MASTER_ID = 103;
defparam axi_monitor_s3.SLAVE_ID = 103;
axi_monitor axi_monitor_s3 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds3_awid         ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awaddr  (ds3_awaddr       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awlen   (ds3_awlen        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awsize  (ds3_awsize       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awburst (ds3_awburst      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awlock  ({1'b0,ds3_awlock}), // () <= ()
	.awcache (ds3_awcache      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awprot  (ds3_awprot       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.awvalid (ds3_awvalid      ), // (axi_monitor_s3,axi_slave3,bench) <= (bmc300)
	.awready (ds3_awready      ), // (axi_monitor_s3,bench,bmc300) <= (axi_slave3)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds3_wid          ), // (axi_monitor_s3,axi_slave3) <= ()
	.wdata   (ds3_wdata        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wstrb   (ds3_wstrb        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wlast   (ds3_wlast        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wvalid  (ds3_wvalid       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.wready  (ds3_wready       ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds3_bid          ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.bresp   (ds3_bresp        ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.bvalid  (ds3_bvalid       ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.bready  (ds3_bready       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds3_arid         ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.araddr  (ds3_araddr       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arlen   (ds3_arlen        ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arsize  (ds3_arsize       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arburst (ds3_arburst      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arlock  ({1'b0,ds3_arlock}), // () <= ()
	.arcache (ds3_arcache      ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arprot  (ds3_arprot       ), // (axi_monitor_s3,axi_slave3) <= (bmc300)
	.arvalid (ds3_arvalid      ), // (axi_monitor_s3,axi_slave3,bench) <= (bmc300)
	.arready (ds3_arready      ), // (axi_monitor_s3,bench,bmc300) <= (axi_slave3)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds3_rid          ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.rdata   (ds3_rdata        ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.rresp   (ds3_rresp        ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.rlast   (ds3_rlast        ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
	.rvalid  (ds3_rvalid       ), // (axi_monitor_s3,bmc300) <= (axi_slave3)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds3_rready       )  // (axi_monitor_s3,axi_slave3) <= (bmc300)
); // end of axi_monitor_s3

`endif // ATCBMC300_SLV3_SUPPORT
`ifdef ATCBMC300_SLV4_SUPPORT
defparam axi_slave4.ADDR_DECODE_WIDTH = `ATCBMC300_SLV4_SIZE+19;
defparam axi_slave4.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave4.AXI4 = 1'b1;
defparam axi_slave4.DATA_WIDTH = DATA_SIZE;
defparam axi_slave4.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave4.MEM_ADDR_WIDTH = `ATCBMC300_SLV4_SIZE+19;
defparam axi_slave4.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave4 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds4_awid         ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awaddr  (ds4_awaddr       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awlen   (ds4_awlen        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awsize  (ds4_awsize       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awburst (ds4_awburst      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awlock  ({1'b0,ds4_awlock}), // () <= ()
	.awcache (ds4_awcache      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awprot  (ds4_awprot       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awvalid (ds4_awvalid      ), // (axi_monitor_s4,axi_slave4,bench) <= (bmc300)
	.awready (ds4_awready      ), // (axi_slave4) => (axi_monitor_s4,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds4_wid          ), // (axi_monitor_s4,axi_slave4) <= ()
	.wdata   (ds4_wdata        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wstrb   (ds4_wstrb        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wlast   (ds4_wlast        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wvalid  (ds4_wvalid       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wready  (ds4_wready       ), // (axi_slave4) => (axi_monitor_s4,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds4_bid          ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.bresp   (ds4_bresp        ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.bvalid  (ds4_bvalid       ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.bready  (ds4_bready       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds4_arid         ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.araddr  (ds4_araddr       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arlen   (ds4_arlen        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arsize  (ds4_arsize       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arburst (ds4_arburst      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arlock  ({1'b0,ds4_arlock}), // () <= ()
	.arcache (ds4_arcache      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arprot  (ds4_arprot       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arvalid (ds4_arvalid      ), // (axi_monitor_s4,axi_slave4,bench) <= (bmc300)
	.arready (ds4_arready      ), // (axi_slave4) => (axi_monitor_s4,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds4_rid          ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.rdata   (ds4_rdata        ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.rresp   (ds4_rresp        ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.rlast   (ds4_rlast        ), // (axi_slave4) => (axi_monitor_s4,bmc300)
	.rvalid  (ds4_rvalid       ), // (axi_slave4) => (axi_monitor_s4,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds4_rready       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave4) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave4

defparam axi_monitor_s4.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s4.AXI4 = 1'b1;
defparam axi_monitor_s4.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s4.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s4.MASTER_ID = 104;
defparam axi_monitor_s4.SLAVE_ID = 104;
axi_monitor axi_monitor_s4 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds4_awid         ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awaddr  (ds4_awaddr       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awlen   (ds4_awlen        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awsize  (ds4_awsize       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awburst (ds4_awburst      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awlock  ({1'b0,ds4_awlock}), // () <= ()
	.awcache (ds4_awcache      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awprot  (ds4_awprot       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.awvalid (ds4_awvalid      ), // (axi_monitor_s4,axi_slave4,bench) <= (bmc300)
	.awready (ds4_awready      ), // (axi_monitor_s4,bench,bmc300) <= (axi_slave4)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds4_wid          ), // (axi_monitor_s4,axi_slave4) <= ()
	.wdata   (ds4_wdata        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wstrb   (ds4_wstrb        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wlast   (ds4_wlast        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wvalid  (ds4_wvalid       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.wready  (ds4_wready       ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds4_bid          ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.bresp   (ds4_bresp        ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.bvalid  (ds4_bvalid       ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.bready  (ds4_bready       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds4_arid         ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.araddr  (ds4_araddr       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arlen   (ds4_arlen        ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arsize  (ds4_arsize       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arburst (ds4_arburst      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arlock  ({1'b0,ds4_arlock}), // () <= ()
	.arcache (ds4_arcache      ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arprot  (ds4_arprot       ), // (axi_monitor_s4,axi_slave4) <= (bmc300)
	.arvalid (ds4_arvalid      ), // (axi_monitor_s4,axi_slave4,bench) <= (bmc300)
	.arready (ds4_arready      ), // (axi_monitor_s4,bench,bmc300) <= (axi_slave4)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds4_rid          ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.rdata   (ds4_rdata        ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.rresp   (ds4_rresp        ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.rlast   (ds4_rlast        ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
	.rvalid  (ds4_rvalid       ), // (axi_monitor_s4,bmc300) <= (axi_slave4)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds4_rready       )  // (axi_monitor_s4,axi_slave4) <= (bmc300)
); // end of axi_monitor_s4

`endif // ATCBMC300_SLV4_SUPPORT
`ifdef ATCBMC300_SLV5_SUPPORT
defparam axi_slave5.ADDR_DECODE_WIDTH = `ATCBMC300_SLV5_SIZE+19;
defparam axi_slave5.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave5.AXI4 = 1'b1;
defparam axi_slave5.DATA_WIDTH = DATA_SIZE;
defparam axi_slave5.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave5.MEM_ADDR_WIDTH = `ATCBMC300_SLV5_SIZE+19;
defparam axi_slave5.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave5 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds5_awid         ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awaddr  (ds5_awaddr       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awlen   (ds5_awlen        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awsize  (ds5_awsize       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awburst (ds5_awburst      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awlock  ({1'b0,ds5_awlock}), // () <= ()
	.awcache (ds5_awcache      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awprot  (ds5_awprot       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awvalid (ds5_awvalid      ), // (axi_monitor_s5,axi_slave5,bench) <= (bmc300)
	.awready (ds5_awready      ), // (axi_slave5) => (axi_monitor_s5,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds5_wid          ), // (axi_monitor_s5,axi_slave5) <= ()
	.wdata   (ds5_wdata        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wstrb   (ds5_wstrb        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wlast   (ds5_wlast        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wvalid  (ds5_wvalid       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wready  (ds5_wready       ), // (axi_slave5) => (axi_monitor_s5,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds5_bid          ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.bresp   (ds5_bresp        ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.bvalid  (ds5_bvalid       ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.bready  (ds5_bready       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds5_arid         ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.araddr  (ds5_araddr       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arlen   (ds5_arlen        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arsize  (ds5_arsize       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arburst (ds5_arburst      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arlock  ({1'b0,ds5_arlock}), // () <= ()
	.arcache (ds5_arcache      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arprot  (ds5_arprot       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arvalid (ds5_arvalid      ), // (axi_monitor_s5,axi_slave5,bench) <= (bmc300)
	.arready (ds5_arready      ), // (axi_slave5) => (axi_monitor_s5,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds5_rid          ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.rdata   (ds5_rdata        ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.rresp   (ds5_rresp        ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.rlast   (ds5_rlast        ), // (axi_slave5) => (axi_monitor_s5,bmc300)
	.rvalid  (ds5_rvalid       ), // (axi_slave5) => (axi_monitor_s5,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds5_rready       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave5) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave5

defparam axi_monitor_s5.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s5.AXI4 = 1'b1;
defparam axi_monitor_s5.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s5.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s5.MASTER_ID = 105;
defparam axi_monitor_s5.SLAVE_ID = 105;
axi_monitor axi_monitor_s5 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds5_awid         ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awaddr  (ds5_awaddr       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awlen   (ds5_awlen        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awsize  (ds5_awsize       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awburst (ds5_awburst      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awlock  ({1'b0,ds5_awlock}), // () <= ()
	.awcache (ds5_awcache      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awprot  (ds5_awprot       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.awvalid (ds5_awvalid      ), // (axi_monitor_s5,axi_slave5,bench) <= (bmc300)
	.awready (ds5_awready      ), // (axi_monitor_s5,bench,bmc300) <= (axi_slave5)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds5_wid          ), // (axi_monitor_s5,axi_slave5) <= ()
	.wdata   (ds5_wdata        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wstrb   (ds5_wstrb        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wlast   (ds5_wlast        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wvalid  (ds5_wvalid       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.wready  (ds5_wready       ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds5_bid          ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.bresp   (ds5_bresp        ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.bvalid  (ds5_bvalid       ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.bready  (ds5_bready       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds5_arid         ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.araddr  (ds5_araddr       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arlen   (ds5_arlen        ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arsize  (ds5_arsize       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arburst (ds5_arburst      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arlock  ({1'b0,ds5_arlock}), // () <= ()
	.arcache (ds5_arcache      ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arprot  (ds5_arprot       ), // (axi_monitor_s5,axi_slave5) <= (bmc300)
	.arvalid (ds5_arvalid      ), // (axi_monitor_s5,axi_slave5,bench) <= (bmc300)
	.arready (ds5_arready      ), // (axi_monitor_s5,bench,bmc300) <= (axi_slave5)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds5_rid          ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.rdata   (ds5_rdata        ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.rresp   (ds5_rresp        ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.rlast   (ds5_rlast        ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
	.rvalid  (ds5_rvalid       ), // (axi_monitor_s5,bmc300) <= (axi_slave5)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds5_rready       )  // (axi_monitor_s5,axi_slave5) <= (bmc300)
); // end of axi_monitor_s5

`endif // ATCBMC300_SLV5_SUPPORT
`ifdef ATCBMC300_SLV6_SUPPORT
defparam axi_slave6.ADDR_DECODE_WIDTH = `ATCBMC300_SLV6_SIZE+19;
defparam axi_slave6.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave6.AXI4 = 1'b1;
defparam axi_slave6.DATA_WIDTH = DATA_SIZE;
defparam axi_slave6.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave6.MEM_ADDR_WIDTH = `ATCBMC300_SLV6_SIZE+19;
defparam axi_slave6.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave6 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds6_awid         ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awaddr  (ds6_awaddr       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awlen   (ds6_awlen        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awsize  (ds6_awsize       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awburst (ds6_awburst      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awlock  ({1'b0,ds6_awlock}), // () <= ()
	.awcache (ds6_awcache      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awprot  (ds6_awprot       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awvalid (ds6_awvalid      ), // (axi_monitor_s6,axi_slave6,bench) <= (bmc300)
	.awready (ds6_awready      ), // (axi_slave6) => (axi_monitor_s6,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds6_wid          ), // (axi_monitor_s6,axi_slave6) <= ()
	.wdata   (ds6_wdata        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wstrb   (ds6_wstrb        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wlast   (ds6_wlast        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wvalid  (ds6_wvalid       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wready  (ds6_wready       ), // (axi_slave6) => (axi_monitor_s6,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds6_bid          ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.bresp   (ds6_bresp        ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.bvalid  (ds6_bvalid       ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.bready  (ds6_bready       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds6_arid         ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.araddr  (ds6_araddr       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arlen   (ds6_arlen        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arsize  (ds6_arsize       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arburst (ds6_arburst      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arlock  ({1'b0,ds6_arlock}), // () <= ()
	.arcache (ds6_arcache      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arprot  (ds6_arprot       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arvalid (ds6_arvalid      ), // (axi_monitor_s6,axi_slave6,bench) <= (bmc300)
	.arready (ds6_arready      ), // (axi_slave6) => (axi_monitor_s6,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds6_rid          ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.rdata   (ds6_rdata        ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.rresp   (ds6_rresp        ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.rlast   (ds6_rlast        ), // (axi_slave6) => (axi_monitor_s6,bmc300)
	.rvalid  (ds6_rvalid       ), // (axi_slave6) => (axi_monitor_s6,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds6_rready       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave6) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave6

defparam axi_monitor_s6.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s6.AXI4 = 1'b1;
defparam axi_monitor_s6.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s6.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s6.MASTER_ID = 106;
defparam axi_monitor_s6.SLAVE_ID = 106;
axi_monitor axi_monitor_s6 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds6_awid         ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awaddr  (ds6_awaddr       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awlen   (ds6_awlen        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awsize  (ds6_awsize       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awburst (ds6_awburst      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awlock  ({1'b0,ds6_awlock}), // () <= ()
	.awcache (ds6_awcache      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awprot  (ds6_awprot       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.awvalid (ds6_awvalid      ), // (axi_monitor_s6,axi_slave6,bench) <= (bmc300)
	.awready (ds6_awready      ), // (axi_monitor_s6,bench,bmc300) <= (axi_slave6)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds6_wid          ), // (axi_monitor_s6,axi_slave6) <= ()
	.wdata   (ds6_wdata        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wstrb   (ds6_wstrb        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wlast   (ds6_wlast        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wvalid  (ds6_wvalid       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.wready  (ds6_wready       ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds6_bid          ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.bresp   (ds6_bresp        ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.bvalid  (ds6_bvalid       ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.bready  (ds6_bready       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds6_arid         ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.araddr  (ds6_araddr       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arlen   (ds6_arlen        ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arsize  (ds6_arsize       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arburst (ds6_arburst      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arlock  ({1'b0,ds6_arlock}), // () <= ()
	.arcache (ds6_arcache      ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arprot  (ds6_arprot       ), // (axi_monitor_s6,axi_slave6) <= (bmc300)
	.arvalid (ds6_arvalid      ), // (axi_monitor_s6,axi_slave6,bench) <= (bmc300)
	.arready (ds6_arready      ), // (axi_monitor_s6,bench,bmc300) <= (axi_slave6)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds6_rid          ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.rdata   (ds6_rdata        ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.rresp   (ds6_rresp        ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.rlast   (ds6_rlast        ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
	.rvalid  (ds6_rvalid       ), // (axi_monitor_s6,bmc300) <= (axi_slave6)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds6_rready       )  // (axi_monitor_s6,axi_slave6) <= (bmc300)
); // end of axi_monitor_s6

`endif // ATCBMC300_SLV6_SUPPORT
`ifdef ATCBMC300_SLV7_SUPPORT
defparam axi_slave7.ADDR_DECODE_WIDTH = `ATCBMC300_SLV7_SIZE+19;
defparam axi_slave7.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave7.AXI4 = 1'b1;
defparam axi_slave7.DATA_WIDTH = DATA_SIZE;
defparam axi_slave7.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave7.MEM_ADDR_WIDTH = `ATCBMC300_SLV7_SIZE+19;
defparam axi_slave7.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave7 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds7_awid         ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awaddr  (ds7_awaddr       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awlen   (ds7_awlen        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awsize  (ds7_awsize       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awburst (ds7_awburst      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awlock  ({1'b0,ds7_awlock}), // () <= ()
	.awcache (ds7_awcache      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awprot  (ds7_awprot       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awvalid (ds7_awvalid      ), // (axi_monitor_s7,axi_slave7,bench) <= (bmc300)
	.awready (ds7_awready      ), // (axi_slave7) => (axi_monitor_s7,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds7_wid          ), // (axi_monitor_s7,axi_slave7) <= ()
	.wdata   (ds7_wdata        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wstrb   (ds7_wstrb        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wlast   (ds7_wlast        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wvalid  (ds7_wvalid       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wready  (ds7_wready       ), // (axi_slave7) => (axi_monitor_s7,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds7_bid          ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.bresp   (ds7_bresp        ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.bvalid  (ds7_bvalid       ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.bready  (ds7_bready       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds7_arid         ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.araddr  (ds7_araddr       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arlen   (ds7_arlen        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arsize  (ds7_arsize       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arburst (ds7_arburst      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arlock  ({1'b0,ds7_arlock}), // () <= ()
	.arcache (ds7_arcache      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arprot  (ds7_arprot       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arvalid (ds7_arvalid      ), // (axi_monitor_s7,axi_slave7,bench) <= (bmc300)
	.arready (ds7_arready      ), // (axi_slave7) => (axi_monitor_s7,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds7_rid          ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.rdata   (ds7_rdata        ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.rresp   (ds7_rresp        ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.rlast   (ds7_rlast        ), // (axi_slave7) => (axi_monitor_s7,bmc300)
	.rvalid  (ds7_rvalid       ), // (axi_slave7) => (axi_monitor_s7,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds7_rready       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave7) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave7

defparam axi_monitor_s7.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s7.AXI4 = 1'b1;
defparam axi_monitor_s7.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s7.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s7.MASTER_ID = 107;
defparam axi_monitor_s7.SLAVE_ID = 107;
axi_monitor axi_monitor_s7 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds7_awid         ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awaddr  (ds7_awaddr       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awlen   (ds7_awlen        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awsize  (ds7_awsize       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awburst (ds7_awburst      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awlock  ({1'b0,ds7_awlock}), // () <= ()
	.awcache (ds7_awcache      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awprot  (ds7_awprot       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.awvalid (ds7_awvalid      ), // (axi_monitor_s7,axi_slave7,bench) <= (bmc300)
	.awready (ds7_awready      ), // (axi_monitor_s7,bench,bmc300) <= (axi_slave7)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds7_wid          ), // (axi_monitor_s7,axi_slave7) <= ()
	.wdata   (ds7_wdata        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wstrb   (ds7_wstrb        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wlast   (ds7_wlast        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wvalid  (ds7_wvalid       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.wready  (ds7_wready       ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds7_bid          ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.bresp   (ds7_bresp        ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.bvalid  (ds7_bvalid       ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.bready  (ds7_bready       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds7_arid         ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.araddr  (ds7_araddr       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arlen   (ds7_arlen        ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arsize  (ds7_arsize       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arburst (ds7_arburst      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arlock  ({1'b0,ds7_arlock}), // () <= ()
	.arcache (ds7_arcache      ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arprot  (ds7_arprot       ), // (axi_monitor_s7,axi_slave7) <= (bmc300)
	.arvalid (ds7_arvalid      ), // (axi_monitor_s7,axi_slave7,bench) <= (bmc300)
	.arready (ds7_arready      ), // (axi_monitor_s7,bench,bmc300) <= (axi_slave7)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds7_rid          ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.rdata   (ds7_rdata        ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.rresp   (ds7_rresp        ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.rlast   (ds7_rlast        ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
	.rvalid  (ds7_rvalid       ), // (axi_monitor_s7,bmc300) <= (axi_slave7)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds7_rready       )  // (axi_monitor_s7,axi_slave7) <= (bmc300)
); // end of axi_monitor_s7

`endif // ATCBMC300_SLV7_SUPPORT
`ifdef ATCBMC300_SLV8_SUPPORT
defparam axi_slave8.ADDR_DECODE_WIDTH = `ATCBMC300_SLV8_SIZE+19;
defparam axi_slave8.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave8.AXI4 = 1'b1;
defparam axi_slave8.DATA_WIDTH = DATA_SIZE;
defparam axi_slave8.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave8.MEM_ADDR_WIDTH = `ATCBMC300_SLV8_SIZE+19;
defparam axi_slave8.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave8 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds8_awid         ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awaddr  (ds8_awaddr       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awlen   (ds8_awlen        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awsize  (ds8_awsize       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awburst (ds8_awburst      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awlock  ({1'b0,ds8_awlock}), // () <= ()
	.awcache (ds8_awcache      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awprot  (ds8_awprot       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awvalid (ds8_awvalid      ), // (axi_monitor_s8,axi_slave8,bench) <= (bmc300)
	.awready (ds8_awready      ), // (axi_slave8) => (axi_monitor_s8,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds8_wid          ), // (axi_monitor_s8,axi_slave8) <= ()
	.wdata   (ds8_wdata        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wstrb   (ds8_wstrb        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wlast   (ds8_wlast        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wvalid  (ds8_wvalid       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wready  (ds8_wready       ), // (axi_slave8) => (axi_monitor_s8,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds8_bid          ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.bresp   (ds8_bresp        ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.bvalid  (ds8_bvalid       ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.bready  (ds8_bready       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds8_arid         ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.araddr  (ds8_araddr       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arlen   (ds8_arlen        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arsize  (ds8_arsize       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arburst (ds8_arburst      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arlock  ({1'b0,ds8_arlock}), // () <= ()
	.arcache (ds8_arcache      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arprot  (ds8_arprot       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arvalid (ds8_arvalid      ), // (axi_monitor_s8,axi_slave8,bench) <= (bmc300)
	.arready (ds8_arready      ), // (axi_slave8) => (axi_monitor_s8,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds8_rid          ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.rdata   (ds8_rdata        ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.rresp   (ds8_rresp        ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.rlast   (ds8_rlast        ), // (axi_slave8) => (axi_monitor_s8,bmc300)
	.rvalid  (ds8_rvalid       ), // (axi_slave8) => (axi_monitor_s8,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds8_rready       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave8) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave8

defparam axi_monitor_s8.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s8.AXI4 = 1'b1;
defparam axi_monitor_s8.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s8.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s8.MASTER_ID = 108;
defparam axi_monitor_s8.SLAVE_ID = 108;
axi_monitor axi_monitor_s8 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds8_awid         ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awaddr  (ds8_awaddr       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awlen   (ds8_awlen        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awsize  (ds8_awsize       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awburst (ds8_awburst      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awlock  ({1'b0,ds8_awlock}), // () <= ()
	.awcache (ds8_awcache      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awprot  (ds8_awprot       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.awvalid (ds8_awvalid      ), // (axi_monitor_s8,axi_slave8,bench) <= (bmc300)
	.awready (ds8_awready      ), // (axi_monitor_s8,bench,bmc300) <= (axi_slave8)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds8_wid          ), // (axi_monitor_s8,axi_slave8) <= ()
	.wdata   (ds8_wdata        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wstrb   (ds8_wstrb        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wlast   (ds8_wlast        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wvalid  (ds8_wvalid       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.wready  (ds8_wready       ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds8_bid          ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.bresp   (ds8_bresp        ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.bvalid  (ds8_bvalid       ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.bready  (ds8_bready       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds8_arid         ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.araddr  (ds8_araddr       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arlen   (ds8_arlen        ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arsize  (ds8_arsize       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arburst (ds8_arburst      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arlock  ({1'b0,ds8_arlock}), // () <= ()
	.arcache (ds8_arcache      ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arprot  (ds8_arprot       ), // (axi_monitor_s8,axi_slave8) <= (bmc300)
	.arvalid (ds8_arvalid      ), // (axi_monitor_s8,axi_slave8,bench) <= (bmc300)
	.arready (ds8_arready      ), // (axi_monitor_s8,bench,bmc300) <= (axi_slave8)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds8_rid          ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.rdata   (ds8_rdata        ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.rresp   (ds8_rresp        ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.rlast   (ds8_rlast        ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
	.rvalid  (ds8_rvalid       ), // (axi_monitor_s8,bmc300) <= (axi_slave8)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds8_rready       )  // (axi_monitor_s8,axi_slave8) <= (bmc300)
); // end of axi_monitor_s8

`endif // ATCBMC300_SLV8_SUPPORT
`ifdef ATCBMC300_SLV9_SUPPORT
defparam axi_slave9.ADDR_DECODE_WIDTH = `ATCBMC300_SLV9_SIZE+19;
defparam axi_slave9.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave9.AXI4 = 1'b1;
defparam axi_slave9.DATA_WIDTH = DATA_SIZE;
defparam axi_slave9.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave9.MEM_ADDR_WIDTH = `ATCBMC300_SLV9_SIZE+19;
defparam axi_slave9.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave9 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds9_awid         ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awaddr  (ds9_awaddr       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awlen   (ds9_awlen        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awsize  (ds9_awsize       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awburst (ds9_awburst      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awlock  ({1'b0,ds9_awlock}), // () <= ()
	.awcache (ds9_awcache      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awprot  (ds9_awprot       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awvalid (ds9_awvalid      ), // (axi_monitor_s9,axi_slave9,bench) <= (bmc300)
	.awready (ds9_awready      ), // (axi_slave9) => (axi_monitor_s9,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds9_wid          ), // (axi_monitor_s9,axi_slave9) <= ()
	.wdata   (ds9_wdata        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wstrb   (ds9_wstrb        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wlast   (ds9_wlast        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wvalid  (ds9_wvalid       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wready  (ds9_wready       ), // (axi_slave9) => (axi_monitor_s9,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds9_bid          ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.bresp   (ds9_bresp        ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.bvalid  (ds9_bvalid       ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.bready  (ds9_bready       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds9_arid         ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.araddr  (ds9_araddr       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arlen   (ds9_arlen        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arsize  (ds9_arsize       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arburst (ds9_arburst      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arlock  ({1'b0,ds9_arlock}), // () <= ()
	.arcache (ds9_arcache      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arprot  (ds9_arprot       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arvalid (ds9_arvalid      ), // (axi_monitor_s9,axi_slave9,bench) <= (bmc300)
	.arready (ds9_arready      ), // (axi_slave9) => (axi_monitor_s9,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds9_rid          ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.rdata   (ds9_rdata        ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.rresp   (ds9_rresp        ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.rlast   (ds9_rlast        ), // (axi_slave9) => (axi_monitor_s9,bmc300)
	.rvalid  (ds9_rvalid       ), // (axi_slave9) => (axi_monitor_s9,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds9_rready       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.csysreq (1'b0             ), // (axi_slave9) <= ()
	.csysack (                 ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                 )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave9

defparam axi_monitor_s9.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s9.AXI4 = 1'b1;
defparam axi_monitor_s9.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s9.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s9.MASTER_ID = 109;
defparam axi_monitor_s9.SLAVE_ID = 109;
axi_monitor axi_monitor_s9 (
	.aclk    (aclk             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn          ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds9_awid         ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awaddr  (ds9_awaddr       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awlen   (ds9_awlen        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awsize  (ds9_awsize       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awburst (ds9_awburst      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awlock  ({1'b0,ds9_awlock}), // () <= ()
	.awcache (ds9_awcache      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awprot  (ds9_awprot       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.awvalid (ds9_awvalid      ), // (axi_monitor_s9,axi_slave9,bench) <= (bmc300)
	.awready (ds9_awready      ), // (axi_monitor_s9,bench,bmc300) <= (axi_slave9)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds9_wid          ), // (axi_monitor_s9,axi_slave9) <= ()
	.wdata   (ds9_wdata        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wstrb   (ds9_wstrb        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wlast   (ds9_wlast        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wvalid  (ds9_wvalid       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.wready  (ds9_wready       ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds9_bid          ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.bresp   (ds9_bresp        ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.bvalid  (ds9_bvalid       ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.bready  (ds9_bready       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds9_arid         ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.araddr  (ds9_araddr       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arlen   (ds9_arlen        ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arsize  (ds9_arsize       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arburst (ds9_arburst      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arlock  ({1'b0,ds9_arlock}), // () <= ()
	.arcache (ds9_arcache      ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arprot  (ds9_arprot       ), // (axi_monitor_s9,axi_slave9) <= (bmc300)
	.arvalid (ds9_arvalid      ), // (axi_monitor_s9,axi_slave9,bench) <= (bmc300)
	.arready (ds9_arready      ), // (axi_monitor_s9,bench,bmc300) <= (axi_slave9)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion         ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser           ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds9_rid          ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.rdata   (ds9_rdata        ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.rresp   (ds9_rresp        ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.rlast   (ds9_rlast        ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
	.rvalid  (ds9_rvalid       ), // (axi_monitor_s9,bmc300) <= (axi_slave9)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser            ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds9_rready       )  // (axi_monitor_s9,axi_slave9) <= (bmc300)
); // end of axi_monitor_s9

`endif // ATCBMC300_SLV9_SUPPORT
`ifdef ATCBMC300_SLV10_SUPPORT
defparam axi_slave10.ADDR_DECODE_WIDTH = `ATCBMC300_SLV10_SIZE+19;
defparam axi_slave10.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave10.AXI4 = 1'b1;
defparam axi_slave10.DATA_WIDTH = DATA_SIZE;
defparam axi_slave10.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave10.MEM_ADDR_WIDTH = `ATCBMC300_SLV10_SIZE+19;
defparam axi_slave10.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave10 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds10_awid         ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awaddr  (ds10_awaddr       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awlen   (ds10_awlen        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awsize  (ds10_awsize       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awburst (ds10_awburst      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awlock  ({1'b0,ds10_awlock}), // () <= ()
	.awcache (ds10_awcache      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awprot  (ds10_awprot       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awvalid (ds10_awvalid      ), // (axi_monitor_s10,axi_slave10,bench) <= (bmc300)
	.awready (ds10_awready      ), // (axi_slave10) => (axi_monitor_s10,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds10_wid          ), // (axi_monitor_s10,axi_slave10) <= ()
	.wdata   (ds10_wdata        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wstrb   (ds10_wstrb        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wlast   (ds10_wlast        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wvalid  (ds10_wvalid       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wready  (ds10_wready       ), // (axi_slave10) => (axi_monitor_s10,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds10_bid          ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.bresp   (ds10_bresp        ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.bvalid  (ds10_bvalid       ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.bready  (ds10_bready       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds10_arid         ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.araddr  (ds10_araddr       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arlen   (ds10_arlen        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arsize  (ds10_arsize       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arburst (ds10_arburst      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arlock  ({1'b0,ds10_arlock}), // () <= ()
	.arcache (ds10_arcache      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arprot  (ds10_arprot       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arvalid (ds10_arvalid      ), // (axi_monitor_s10,axi_slave10,bench) <= (bmc300)
	.arready (ds10_arready      ), // (axi_slave10) => (axi_monitor_s10,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds10_rid          ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.rdata   (ds10_rdata        ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.rresp   (ds10_rresp        ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.rlast   (ds10_rlast        ), // (axi_slave10) => (axi_monitor_s10,bmc300)
	.rvalid  (ds10_rvalid       ), // (axi_slave10) => (axi_monitor_s10,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds10_rready       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave10) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave10

defparam axi_monitor_s10.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s10.AXI4 = 1'b1;
defparam axi_monitor_s10.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s10.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s10.MASTER_ID = 110;
defparam axi_monitor_s10.SLAVE_ID = 110;
axi_monitor axi_monitor_s10 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds10_awid         ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awaddr  (ds10_awaddr       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awlen   (ds10_awlen        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awsize  (ds10_awsize       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awburst (ds10_awburst      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awlock  ({1'b0,ds10_awlock}), // () <= ()
	.awcache (ds10_awcache      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awprot  (ds10_awprot       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.awvalid (ds10_awvalid      ), // (axi_monitor_s10,axi_slave10,bench) <= (bmc300)
	.awready (ds10_awready      ), // (axi_monitor_s10,bench,bmc300) <= (axi_slave10)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds10_wid          ), // (axi_monitor_s10,axi_slave10) <= ()
	.wdata   (ds10_wdata        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wstrb   (ds10_wstrb        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wlast   (ds10_wlast        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wvalid  (ds10_wvalid       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.wready  (ds10_wready       ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds10_bid          ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.bresp   (ds10_bresp        ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.bvalid  (ds10_bvalid       ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.bready  (ds10_bready       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds10_arid         ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.araddr  (ds10_araddr       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arlen   (ds10_arlen        ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arsize  (ds10_arsize       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arburst (ds10_arburst      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arlock  ({1'b0,ds10_arlock}), // () <= ()
	.arcache (ds10_arcache      ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arprot  (ds10_arprot       ), // (axi_monitor_s10,axi_slave10) <= (bmc300)
	.arvalid (ds10_arvalid      ), // (axi_monitor_s10,axi_slave10,bench) <= (bmc300)
	.arready (ds10_arready      ), // (axi_monitor_s10,bench,bmc300) <= (axi_slave10)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds10_rid          ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.rdata   (ds10_rdata        ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.rresp   (ds10_rresp        ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.rlast   (ds10_rlast        ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
	.rvalid  (ds10_rvalid       ), // (axi_monitor_s10,bmc300) <= (axi_slave10)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds10_rready       )  // (axi_monitor_s10,axi_slave10) <= (bmc300)
); // end of axi_monitor_s10

`endif // ATCBMC300_SLV10_SUPPORT
`ifdef ATCBMC300_SLV11_SUPPORT
defparam axi_slave11.ADDR_DECODE_WIDTH = `ATCBMC300_SLV11_SIZE+19;
defparam axi_slave11.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave11.AXI4 = 1'b1;
defparam axi_slave11.DATA_WIDTH = DATA_SIZE;
defparam axi_slave11.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave11.MEM_ADDR_WIDTH = `ATCBMC300_SLV11_SIZE+19;
defparam axi_slave11.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave11 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds11_awid         ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awaddr  (ds11_awaddr       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awlen   (ds11_awlen        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awsize  (ds11_awsize       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awburst (ds11_awburst      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awlock  ({1'b0,ds11_awlock}), // () <= ()
	.awcache (ds11_awcache      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awprot  (ds11_awprot       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awvalid (ds11_awvalid      ), // (axi_monitor_s11,axi_slave11,bench) <= (bmc300)
	.awready (ds11_awready      ), // (axi_slave11) => (axi_monitor_s11,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds11_wid          ), // (axi_monitor_s11,axi_slave11) <= ()
	.wdata   (ds11_wdata        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wstrb   (ds11_wstrb        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wlast   (ds11_wlast        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wvalid  (ds11_wvalid       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wready  (ds11_wready       ), // (axi_slave11) => (axi_monitor_s11,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds11_bid          ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.bresp   (ds11_bresp        ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.bvalid  (ds11_bvalid       ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.bready  (ds11_bready       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds11_arid         ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.araddr  (ds11_araddr       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arlen   (ds11_arlen        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arsize  (ds11_arsize       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arburst (ds11_arburst      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arlock  ({1'b0,ds11_arlock}), // () <= ()
	.arcache (ds11_arcache      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arprot  (ds11_arprot       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arvalid (ds11_arvalid      ), // (axi_monitor_s11,axi_slave11,bench) <= (bmc300)
	.arready (ds11_arready      ), // (axi_slave11) => (axi_monitor_s11,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds11_rid          ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.rdata   (ds11_rdata        ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.rresp   (ds11_rresp        ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.rlast   (ds11_rlast        ), // (axi_slave11) => (axi_monitor_s11,bmc300)
	.rvalid  (ds11_rvalid       ), // (axi_slave11) => (axi_monitor_s11,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds11_rready       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave11) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave11

defparam axi_monitor_s11.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s11.AXI4 = 1'b1;
defparam axi_monitor_s11.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s11.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s11.MASTER_ID = 111;
defparam axi_monitor_s11.SLAVE_ID = 111;
axi_monitor axi_monitor_s11 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds11_awid         ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awaddr  (ds11_awaddr       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awlen   (ds11_awlen        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awsize  (ds11_awsize       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awburst (ds11_awburst      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awlock  ({1'b0,ds11_awlock}), // () <= ()
	.awcache (ds11_awcache      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awprot  (ds11_awprot       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.awvalid (ds11_awvalid      ), // (axi_monitor_s11,axi_slave11,bench) <= (bmc300)
	.awready (ds11_awready      ), // (axi_monitor_s11,bench,bmc300) <= (axi_slave11)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds11_wid          ), // (axi_monitor_s11,axi_slave11) <= ()
	.wdata   (ds11_wdata        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wstrb   (ds11_wstrb        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wlast   (ds11_wlast        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wvalid  (ds11_wvalid       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.wready  (ds11_wready       ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds11_bid          ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.bresp   (ds11_bresp        ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.bvalid  (ds11_bvalid       ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.bready  (ds11_bready       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds11_arid         ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.araddr  (ds11_araddr       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arlen   (ds11_arlen        ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arsize  (ds11_arsize       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arburst (ds11_arburst      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arlock  ({1'b0,ds11_arlock}), // () <= ()
	.arcache (ds11_arcache      ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arprot  (ds11_arprot       ), // (axi_monitor_s11,axi_slave11) <= (bmc300)
	.arvalid (ds11_arvalid      ), // (axi_monitor_s11,axi_slave11,bench) <= (bmc300)
	.arready (ds11_arready      ), // (axi_monitor_s11,bench,bmc300) <= (axi_slave11)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds11_rid          ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.rdata   (ds11_rdata        ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.rresp   (ds11_rresp        ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.rlast   (ds11_rlast        ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
	.rvalid  (ds11_rvalid       ), // (axi_monitor_s11,bmc300) <= (axi_slave11)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds11_rready       )  // (axi_monitor_s11,axi_slave11) <= (bmc300)
); // end of axi_monitor_s11

`endif // ATCBMC300_SLV11_SUPPORT
`ifdef ATCBMC300_SLV12_SUPPORT
defparam axi_slave12.ADDR_DECODE_WIDTH = `ATCBMC300_SLV12_SIZE+19;
defparam axi_slave12.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave12.AXI4 = 1'b1;
defparam axi_slave12.DATA_WIDTH = DATA_SIZE;
defparam axi_slave12.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave12.MEM_ADDR_WIDTH = `ATCBMC300_SLV12_SIZE+19;
defparam axi_slave12.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave12 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds12_awid         ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awaddr  (ds12_awaddr       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awlen   (ds12_awlen        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awsize  (ds12_awsize       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awburst (ds12_awburst      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awlock  ({1'b0,ds12_awlock}), // () <= ()
	.awcache (ds12_awcache      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awprot  (ds12_awprot       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awvalid (ds12_awvalid      ), // (axi_monitor_s12,axi_slave12,bench) <= (bmc300)
	.awready (ds12_awready      ), // (axi_slave12) => (axi_monitor_s12,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds12_wid          ), // (axi_monitor_s12,axi_slave12) <= ()
	.wdata   (ds12_wdata        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wstrb   (ds12_wstrb        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wlast   (ds12_wlast        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wvalid  (ds12_wvalid       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wready  (ds12_wready       ), // (axi_slave12) => (axi_monitor_s12,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds12_bid          ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.bresp   (ds12_bresp        ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.bvalid  (ds12_bvalid       ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.bready  (ds12_bready       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds12_arid         ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.araddr  (ds12_araddr       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arlen   (ds12_arlen        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arsize  (ds12_arsize       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arburst (ds12_arburst      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arlock  ({1'b0,ds12_arlock}), // () <= ()
	.arcache (ds12_arcache      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arprot  (ds12_arprot       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arvalid (ds12_arvalid      ), // (axi_monitor_s12,axi_slave12,bench) <= (bmc300)
	.arready (ds12_arready      ), // (axi_slave12) => (axi_monitor_s12,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds12_rid          ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.rdata   (ds12_rdata        ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.rresp   (ds12_rresp        ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.rlast   (ds12_rlast        ), // (axi_slave12) => (axi_monitor_s12,bmc300)
	.rvalid  (ds12_rvalid       ), // (axi_slave12) => (axi_monitor_s12,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds12_rready       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave12) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave12

defparam axi_monitor_s12.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s12.AXI4 = 1'b1;
defparam axi_monitor_s12.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s12.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s12.MASTER_ID = 112;
defparam axi_monitor_s12.SLAVE_ID = 112;
axi_monitor axi_monitor_s12 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds12_awid         ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awaddr  (ds12_awaddr       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awlen   (ds12_awlen        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awsize  (ds12_awsize       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awburst (ds12_awburst      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awlock  ({1'b0,ds12_awlock}), // () <= ()
	.awcache (ds12_awcache      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awprot  (ds12_awprot       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.awvalid (ds12_awvalid      ), // (axi_monitor_s12,axi_slave12,bench) <= (bmc300)
	.awready (ds12_awready      ), // (axi_monitor_s12,bench,bmc300) <= (axi_slave12)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds12_wid          ), // (axi_monitor_s12,axi_slave12) <= ()
	.wdata   (ds12_wdata        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wstrb   (ds12_wstrb        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wlast   (ds12_wlast        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wvalid  (ds12_wvalid       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.wready  (ds12_wready       ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds12_bid          ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.bresp   (ds12_bresp        ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.bvalid  (ds12_bvalid       ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.bready  (ds12_bready       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds12_arid         ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.araddr  (ds12_araddr       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arlen   (ds12_arlen        ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arsize  (ds12_arsize       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arburst (ds12_arburst      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arlock  ({1'b0,ds12_arlock}), // () <= ()
	.arcache (ds12_arcache      ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arprot  (ds12_arprot       ), // (axi_monitor_s12,axi_slave12) <= (bmc300)
	.arvalid (ds12_arvalid      ), // (axi_monitor_s12,axi_slave12,bench) <= (bmc300)
	.arready (ds12_arready      ), // (axi_monitor_s12,bench,bmc300) <= (axi_slave12)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds12_rid          ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.rdata   (ds12_rdata        ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.rresp   (ds12_rresp        ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.rlast   (ds12_rlast        ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
	.rvalid  (ds12_rvalid       ), // (axi_monitor_s12,bmc300) <= (axi_slave12)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds12_rready       )  // (axi_monitor_s12,axi_slave12) <= (bmc300)
); // end of axi_monitor_s12

`endif // ATCBMC300_SLV12_SUPPORT
`ifdef ATCBMC300_SLV13_SUPPORT
defparam axi_slave13.ADDR_DECODE_WIDTH = `ATCBMC300_SLV13_SIZE+19;
defparam axi_slave13.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave13.AXI4 = 1'b1;
defparam axi_slave13.DATA_WIDTH = DATA_SIZE;
defparam axi_slave13.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave13.MEM_ADDR_WIDTH = `ATCBMC300_SLV13_SIZE+19;
defparam axi_slave13.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave13 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds13_awid         ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awaddr  (ds13_awaddr       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awlen   (ds13_awlen        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awsize  (ds13_awsize       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awburst (ds13_awburst      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awlock  ({1'b0,ds13_awlock}), // () <= ()
	.awcache (ds13_awcache      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awprot  (ds13_awprot       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awvalid (ds13_awvalid      ), // (axi_monitor_s13,axi_slave13,bench) <= (bmc300)
	.awready (ds13_awready      ), // (axi_slave13) => (axi_monitor_s13,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds13_wid          ), // (axi_monitor_s13,axi_slave13) <= ()
	.wdata   (ds13_wdata        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wstrb   (ds13_wstrb        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wlast   (ds13_wlast        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wvalid  (ds13_wvalid       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wready  (ds13_wready       ), // (axi_slave13) => (axi_monitor_s13,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds13_bid          ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.bresp   (ds13_bresp        ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.bvalid  (ds13_bvalid       ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.bready  (ds13_bready       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds13_arid         ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.araddr  (ds13_araddr       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arlen   (ds13_arlen        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arsize  (ds13_arsize       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arburst (ds13_arburst      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arlock  ({1'b0,ds13_arlock}), // () <= ()
	.arcache (ds13_arcache      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arprot  (ds13_arprot       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arvalid (ds13_arvalid      ), // (axi_monitor_s13,axi_slave13,bench) <= (bmc300)
	.arready (ds13_arready      ), // (axi_slave13) => (axi_monitor_s13,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds13_rid          ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.rdata   (ds13_rdata        ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.rresp   (ds13_rresp        ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.rlast   (ds13_rlast        ), // (axi_slave13) => (axi_monitor_s13,bmc300)
	.rvalid  (ds13_rvalid       ), // (axi_slave13) => (axi_monitor_s13,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds13_rready       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave13) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave13

defparam axi_monitor_s13.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s13.AXI4 = 1'b1;
defparam axi_monitor_s13.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s13.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s13.MASTER_ID = 113;
defparam axi_monitor_s13.SLAVE_ID = 113;
axi_monitor axi_monitor_s13 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds13_awid         ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awaddr  (ds13_awaddr       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awlen   (ds13_awlen        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awsize  (ds13_awsize       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awburst (ds13_awburst      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awlock  ({1'b0,ds13_awlock}), // () <= ()
	.awcache (ds13_awcache      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awprot  (ds13_awprot       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.awvalid (ds13_awvalid      ), // (axi_monitor_s13,axi_slave13,bench) <= (bmc300)
	.awready (ds13_awready      ), // (axi_monitor_s13,bench,bmc300) <= (axi_slave13)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds13_wid          ), // (axi_monitor_s13,axi_slave13) <= ()
	.wdata   (ds13_wdata        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wstrb   (ds13_wstrb        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wlast   (ds13_wlast        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wvalid  (ds13_wvalid       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.wready  (ds13_wready       ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds13_bid          ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.bresp   (ds13_bresp        ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.bvalid  (ds13_bvalid       ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.bready  (ds13_bready       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds13_arid         ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.araddr  (ds13_araddr       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arlen   (ds13_arlen        ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arsize  (ds13_arsize       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arburst (ds13_arburst      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arlock  ({1'b0,ds13_arlock}), // () <= ()
	.arcache (ds13_arcache      ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arprot  (ds13_arprot       ), // (axi_monitor_s13,axi_slave13) <= (bmc300)
	.arvalid (ds13_arvalid      ), // (axi_monitor_s13,axi_slave13,bench) <= (bmc300)
	.arready (ds13_arready      ), // (axi_monitor_s13,bench,bmc300) <= (axi_slave13)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds13_rid          ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.rdata   (ds13_rdata        ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.rresp   (ds13_rresp        ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.rlast   (ds13_rlast        ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
	.rvalid  (ds13_rvalid       ), // (axi_monitor_s13,bmc300) <= (axi_slave13)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds13_rready       )  // (axi_monitor_s13,axi_slave13) <= (bmc300)
); // end of axi_monitor_s13

`endif // ATCBMC300_SLV13_SUPPORT
`ifdef ATCBMC300_SLV14_SUPPORT
defparam axi_slave14.ADDR_DECODE_WIDTH = `ATCBMC300_SLV14_SIZE+19;
defparam axi_slave14.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave14.AXI4 = 1'b1;
defparam axi_slave14.DATA_WIDTH = DATA_SIZE;
defparam axi_slave14.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave14.MEM_ADDR_WIDTH = `ATCBMC300_SLV14_SIZE+19;
defparam axi_slave14.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave14 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds14_awid         ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awaddr  (ds14_awaddr       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awlen   (ds14_awlen        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awsize  (ds14_awsize       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awburst (ds14_awburst      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awlock  ({1'b0,ds14_awlock}), // () <= ()
	.awcache (ds14_awcache      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awprot  (ds14_awprot       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awvalid (ds14_awvalid      ), // (axi_monitor_s14,axi_slave14,bench) <= (bmc300)
	.awready (ds14_awready      ), // (axi_slave14) => (axi_monitor_s14,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds14_wid          ), // (axi_monitor_s14,axi_slave14) <= ()
	.wdata   (ds14_wdata        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wstrb   (ds14_wstrb        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wlast   (ds14_wlast        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wvalid  (ds14_wvalid       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wready  (ds14_wready       ), // (axi_slave14) => (axi_monitor_s14,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds14_bid          ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.bresp   (ds14_bresp        ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.bvalid  (ds14_bvalid       ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.bready  (ds14_bready       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds14_arid         ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.araddr  (ds14_araddr       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arlen   (ds14_arlen        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arsize  (ds14_arsize       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arburst (ds14_arburst      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arlock  ({1'b0,ds14_arlock}), // () <= ()
	.arcache (ds14_arcache      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arprot  (ds14_arprot       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arvalid (ds14_arvalid      ), // (axi_monitor_s14,axi_slave14,bench) <= (bmc300)
	.arready (ds14_arready      ), // (axi_slave14) => (axi_monitor_s14,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds14_rid          ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.rdata   (ds14_rdata        ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.rresp   (ds14_rresp        ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.rlast   (ds14_rlast        ), // (axi_slave14) => (axi_monitor_s14,bmc300)
	.rvalid  (ds14_rvalid       ), // (axi_slave14) => (axi_monitor_s14,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds14_rready       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave14) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave14

defparam axi_monitor_s14.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s14.AXI4 = 1'b1;
defparam axi_monitor_s14.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s14.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s14.MASTER_ID = 114;
defparam axi_monitor_s14.SLAVE_ID = 114;
axi_monitor axi_monitor_s14 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds14_awid         ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awaddr  (ds14_awaddr       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awlen   (ds14_awlen        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awsize  (ds14_awsize       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awburst (ds14_awburst      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awlock  ({1'b0,ds14_awlock}), // () <= ()
	.awcache (ds14_awcache      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awprot  (ds14_awprot       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.awvalid (ds14_awvalid      ), // (axi_monitor_s14,axi_slave14,bench) <= (bmc300)
	.awready (ds14_awready      ), // (axi_monitor_s14,bench,bmc300) <= (axi_slave14)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds14_wid          ), // (axi_monitor_s14,axi_slave14) <= ()
	.wdata   (ds14_wdata        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wstrb   (ds14_wstrb        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wlast   (ds14_wlast        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wvalid  (ds14_wvalid       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.wready  (ds14_wready       ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds14_bid          ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.bresp   (ds14_bresp        ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.bvalid  (ds14_bvalid       ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.bready  (ds14_bready       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds14_arid         ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.araddr  (ds14_araddr       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arlen   (ds14_arlen        ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arsize  (ds14_arsize       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arburst (ds14_arburst      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arlock  ({1'b0,ds14_arlock}), // () <= ()
	.arcache (ds14_arcache      ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arprot  (ds14_arprot       ), // (axi_monitor_s14,axi_slave14) <= (bmc300)
	.arvalid (ds14_arvalid      ), // (axi_monitor_s14,axi_slave14,bench) <= (bmc300)
	.arready (ds14_arready      ), // (axi_monitor_s14,bench,bmc300) <= (axi_slave14)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds14_rid          ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.rdata   (ds14_rdata        ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.rresp   (ds14_rresp        ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.rlast   (ds14_rlast        ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
	.rvalid  (ds14_rvalid       ), // (axi_monitor_s14,bmc300) <= (axi_slave14)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds14_rready       )  // (axi_monitor_s14,axi_slave14) <= (bmc300)
); // end of axi_monitor_s14

`endif // ATCBMC300_SLV14_SUPPORT
`ifdef ATCBMC300_SLV15_SUPPORT
defparam axi_slave15.ADDR_DECODE_WIDTH = `ATCBMC300_SLV15_SIZE+19;
defparam axi_slave15.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave15.AXI4 = 1'b1;
defparam axi_slave15.DATA_WIDTH = DATA_SIZE;
defparam axi_slave15.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave15.MEM_ADDR_WIDTH = `ATCBMC300_SLV15_SIZE+19;
defparam axi_slave15.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave15 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds15_awid         ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awaddr  (ds15_awaddr       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awlen   (ds15_awlen        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awsize  (ds15_awsize       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awburst (ds15_awburst      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awlock  ({1'b0,ds15_awlock}), // () <= ()
	.awcache (ds15_awcache      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awprot  (ds15_awprot       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awvalid (ds15_awvalid      ), // (axi_monitor_s15,axi_slave15,bench) <= (bmc300)
	.awready (ds15_awready      ), // (axi_slave15) => (axi_monitor_s15,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds15_wid          ), // (axi_monitor_s15,axi_slave15) <= ()
	.wdata   (ds15_wdata        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wstrb   (ds15_wstrb        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wlast   (ds15_wlast        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wvalid  (ds15_wvalid       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wready  (ds15_wready       ), // (axi_slave15) => (axi_monitor_s15,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds15_bid          ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.bresp   (ds15_bresp        ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.bvalid  (ds15_bvalid       ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.bready  (ds15_bready       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds15_arid         ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.araddr  (ds15_araddr       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arlen   (ds15_arlen        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arsize  (ds15_arsize       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arburst (ds15_arburst      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arlock  ({1'b0,ds15_arlock}), // () <= ()
	.arcache (ds15_arcache      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arprot  (ds15_arprot       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arvalid (ds15_arvalid      ), // (axi_monitor_s15,axi_slave15,bench) <= (bmc300)
	.arready (ds15_arready      ), // (axi_slave15) => (axi_monitor_s15,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds15_rid          ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.rdata   (ds15_rdata        ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.rresp   (ds15_rresp        ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.rlast   (ds15_rlast        ), // (axi_slave15) => (axi_monitor_s15,bmc300)
	.rvalid  (ds15_rvalid       ), // (axi_slave15) => (axi_monitor_s15,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds15_rready       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave15) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave15

defparam axi_monitor_s15.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s15.AXI4 = 1'b1;
defparam axi_monitor_s15.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s15.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s15.MASTER_ID = 115;
defparam axi_monitor_s15.SLAVE_ID = 115;
axi_monitor axi_monitor_s15 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds15_awid         ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awaddr  (ds15_awaddr       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awlen   (ds15_awlen        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awsize  (ds15_awsize       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awburst (ds15_awburst      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awlock  ({1'b0,ds15_awlock}), // () <= ()
	.awcache (ds15_awcache      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awprot  (ds15_awprot       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.awvalid (ds15_awvalid      ), // (axi_monitor_s15,axi_slave15,bench) <= (bmc300)
	.awready (ds15_awready      ), // (axi_monitor_s15,bench,bmc300) <= (axi_slave15)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds15_wid          ), // (axi_monitor_s15,axi_slave15) <= ()
	.wdata   (ds15_wdata        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wstrb   (ds15_wstrb        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wlast   (ds15_wlast        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wvalid  (ds15_wvalid       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.wready  (ds15_wready       ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds15_bid          ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.bresp   (ds15_bresp        ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.bvalid  (ds15_bvalid       ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.bready  (ds15_bready       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds15_arid         ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.araddr  (ds15_araddr       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arlen   (ds15_arlen        ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arsize  (ds15_arsize       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arburst (ds15_arburst      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arlock  ({1'b0,ds15_arlock}), // () <= ()
	.arcache (ds15_arcache      ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arprot  (ds15_arprot       ), // (axi_monitor_s15,axi_slave15) <= (bmc300)
	.arvalid (ds15_arvalid      ), // (axi_monitor_s15,axi_slave15,bench) <= (bmc300)
	.arready (ds15_arready      ), // (axi_monitor_s15,bench,bmc300) <= (axi_slave15)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds15_rid          ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.rdata   (ds15_rdata        ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.rresp   (ds15_rresp        ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.rlast   (ds15_rlast        ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
	.rvalid  (ds15_rvalid       ), // (axi_monitor_s15,bmc300) <= (axi_slave15)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds15_rready       )  // (axi_monitor_s15,axi_slave15) <= (bmc300)
); // end of axi_monitor_s15

`endif // ATCBMC300_SLV15_SUPPORT
`ifdef ATCBMC300_SLV16_SUPPORT
defparam axi_slave16.ADDR_DECODE_WIDTH = `ATCBMC300_SLV16_SIZE+19;
defparam axi_slave16.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave16.AXI4 = 1'b1;
defparam axi_slave16.DATA_WIDTH = DATA_SIZE;
defparam axi_slave16.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave16.MEM_ADDR_WIDTH = `ATCBMC300_SLV16_SIZE+19;
defparam axi_slave16.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave16 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds16_awid         ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awaddr  (ds16_awaddr       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awlen   (ds16_awlen        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awsize  (ds16_awsize       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awburst (ds16_awburst      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awlock  ({1'b0,ds16_awlock}), // () <= ()
	.awcache (ds16_awcache      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awprot  (ds16_awprot       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awvalid (ds16_awvalid      ), // (axi_monitor_s16,axi_slave16,bench) <= (bmc300)
	.awready (ds16_awready      ), // (axi_slave16) => (axi_monitor_s16,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds16_wid          ), // (axi_monitor_s16,axi_slave16) <= ()
	.wdata   (ds16_wdata        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wstrb   (ds16_wstrb        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wlast   (ds16_wlast        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wvalid  (ds16_wvalid       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wready  (ds16_wready       ), // (axi_slave16) => (axi_monitor_s16,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds16_bid          ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.bresp   (ds16_bresp        ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.bvalid  (ds16_bvalid       ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.bready  (ds16_bready       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds16_arid         ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.araddr  (ds16_araddr       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arlen   (ds16_arlen        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arsize  (ds16_arsize       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arburst (ds16_arburst      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arlock  ({1'b0,ds16_arlock}), // () <= ()
	.arcache (ds16_arcache      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arprot  (ds16_arprot       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arvalid (ds16_arvalid      ), // (axi_monitor_s16,axi_slave16,bench) <= (bmc300)
	.arready (ds16_arready      ), // (axi_slave16) => (axi_monitor_s16,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds16_rid          ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.rdata   (ds16_rdata        ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.rresp   (ds16_rresp        ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.rlast   (ds16_rlast        ), // (axi_slave16) => (axi_monitor_s16,bmc300)
	.rvalid  (ds16_rvalid       ), // (axi_slave16) => (axi_monitor_s16,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds16_rready       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave16) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave16

defparam axi_monitor_s16.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s16.AXI4 = 1'b1;
defparam axi_monitor_s16.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s16.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s16.MASTER_ID = 116;
defparam axi_monitor_s16.SLAVE_ID = 116;
axi_monitor axi_monitor_s16 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds16_awid         ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awaddr  (ds16_awaddr       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awlen   (ds16_awlen        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awsize  (ds16_awsize       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awburst (ds16_awburst      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awlock  ({1'b0,ds16_awlock}), // () <= ()
	.awcache (ds16_awcache      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awprot  (ds16_awprot       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.awvalid (ds16_awvalid      ), // (axi_monitor_s16,axi_slave16,bench) <= (bmc300)
	.awready (ds16_awready      ), // (axi_monitor_s16,bench,bmc300) <= (axi_slave16)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds16_wid          ), // (axi_monitor_s16,axi_slave16) <= ()
	.wdata   (ds16_wdata        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wstrb   (ds16_wstrb        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wlast   (ds16_wlast        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wvalid  (ds16_wvalid       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.wready  (ds16_wready       ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds16_bid          ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.bresp   (ds16_bresp        ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.bvalid  (ds16_bvalid       ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.bready  (ds16_bready       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds16_arid         ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.araddr  (ds16_araddr       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arlen   (ds16_arlen        ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arsize  (ds16_arsize       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arburst (ds16_arburst      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arlock  ({1'b0,ds16_arlock}), // () <= ()
	.arcache (ds16_arcache      ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arprot  (ds16_arprot       ), // (axi_monitor_s16,axi_slave16) <= (bmc300)
	.arvalid (ds16_arvalid      ), // (axi_monitor_s16,axi_slave16,bench) <= (bmc300)
	.arready (ds16_arready      ), // (axi_monitor_s16,bench,bmc300) <= (axi_slave16)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds16_rid          ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.rdata   (ds16_rdata        ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.rresp   (ds16_rresp        ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.rlast   (ds16_rlast        ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
	.rvalid  (ds16_rvalid       ), // (axi_monitor_s16,bmc300) <= (axi_slave16)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds16_rready       )  // (axi_monitor_s16,axi_slave16) <= (bmc300)
); // end of axi_monitor_s16

`endif // ATCBMC300_SLV16_SUPPORT
`ifdef ATCBMC300_SLV17_SUPPORT
defparam axi_slave17.ADDR_DECODE_WIDTH = `ATCBMC300_SLV17_SIZE+19;
defparam axi_slave17.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave17.AXI4 = 1'b1;
defparam axi_slave17.DATA_WIDTH = DATA_SIZE;
defparam axi_slave17.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave17.MEM_ADDR_WIDTH = `ATCBMC300_SLV17_SIZE+19;
defparam axi_slave17.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave17 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds17_awid         ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awaddr  (ds17_awaddr       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awlen   (ds17_awlen        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awsize  (ds17_awsize       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awburst (ds17_awburst      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awlock  ({1'b0,ds17_awlock}), // () <= ()
	.awcache (ds17_awcache      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awprot  (ds17_awprot       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awvalid (ds17_awvalid      ), // (axi_monitor_s17,axi_slave17,bench) <= (bmc300)
	.awready (ds17_awready      ), // (axi_slave17) => (axi_monitor_s17,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds17_wid          ), // (axi_monitor_s17,axi_slave17) <= ()
	.wdata   (ds17_wdata        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wstrb   (ds17_wstrb        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wlast   (ds17_wlast        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wvalid  (ds17_wvalid       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wready  (ds17_wready       ), // (axi_slave17) => (axi_monitor_s17,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds17_bid          ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.bresp   (ds17_bresp        ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.bvalid  (ds17_bvalid       ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.bready  (ds17_bready       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds17_arid         ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.araddr  (ds17_araddr       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arlen   (ds17_arlen        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arsize  (ds17_arsize       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arburst (ds17_arburst      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arlock  ({1'b0,ds17_arlock}), // () <= ()
	.arcache (ds17_arcache      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arprot  (ds17_arprot       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arvalid (ds17_arvalid      ), // (axi_monitor_s17,axi_slave17,bench) <= (bmc300)
	.arready (ds17_arready      ), // (axi_slave17) => (axi_monitor_s17,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds17_rid          ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.rdata   (ds17_rdata        ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.rresp   (ds17_rresp        ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.rlast   (ds17_rlast        ), // (axi_slave17) => (axi_monitor_s17,bmc300)
	.rvalid  (ds17_rvalid       ), // (axi_slave17) => (axi_monitor_s17,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds17_rready       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave17) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave17

defparam axi_monitor_s17.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s17.AXI4 = 1'b1;
defparam axi_monitor_s17.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s17.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s17.MASTER_ID = 117;
defparam axi_monitor_s17.SLAVE_ID = 117;
axi_monitor axi_monitor_s17 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds17_awid         ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awaddr  (ds17_awaddr       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awlen   (ds17_awlen        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awsize  (ds17_awsize       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awburst (ds17_awburst      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awlock  ({1'b0,ds17_awlock}), // () <= ()
	.awcache (ds17_awcache      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awprot  (ds17_awprot       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.awvalid (ds17_awvalid      ), // (axi_monitor_s17,axi_slave17,bench) <= (bmc300)
	.awready (ds17_awready      ), // (axi_monitor_s17,bench,bmc300) <= (axi_slave17)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds17_wid          ), // (axi_monitor_s17,axi_slave17) <= ()
	.wdata   (ds17_wdata        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wstrb   (ds17_wstrb        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wlast   (ds17_wlast        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wvalid  (ds17_wvalid       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.wready  (ds17_wready       ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds17_bid          ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.bresp   (ds17_bresp        ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.bvalid  (ds17_bvalid       ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.bready  (ds17_bready       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds17_arid         ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.araddr  (ds17_araddr       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arlen   (ds17_arlen        ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arsize  (ds17_arsize       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arburst (ds17_arburst      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arlock  ({1'b0,ds17_arlock}), // () <= ()
	.arcache (ds17_arcache      ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arprot  (ds17_arprot       ), // (axi_monitor_s17,axi_slave17) <= (bmc300)
	.arvalid (ds17_arvalid      ), // (axi_monitor_s17,axi_slave17,bench) <= (bmc300)
	.arready (ds17_arready      ), // (axi_monitor_s17,bench,bmc300) <= (axi_slave17)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds17_rid          ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.rdata   (ds17_rdata        ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.rresp   (ds17_rresp        ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.rlast   (ds17_rlast        ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
	.rvalid  (ds17_rvalid       ), // (axi_monitor_s17,bmc300) <= (axi_slave17)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds17_rready       )  // (axi_monitor_s17,axi_slave17) <= (bmc300)
); // end of axi_monitor_s17

`endif // ATCBMC300_SLV17_SUPPORT
`ifdef ATCBMC300_SLV18_SUPPORT
defparam axi_slave18.ADDR_DECODE_WIDTH = `ATCBMC300_SLV18_SIZE+19;
defparam axi_slave18.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave18.AXI4 = 1'b1;
defparam axi_slave18.DATA_WIDTH = DATA_SIZE;
defparam axi_slave18.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave18.MEM_ADDR_WIDTH = `ATCBMC300_SLV18_SIZE+19;
defparam axi_slave18.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave18 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds18_awid         ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awaddr  (ds18_awaddr       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awlen   (ds18_awlen        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awsize  (ds18_awsize       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awburst (ds18_awburst      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awlock  ({1'b0,ds18_awlock}), // () <= ()
	.awcache (ds18_awcache      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awprot  (ds18_awprot       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awvalid (ds18_awvalid      ), // (axi_monitor_s18,axi_slave18,bench) <= (bmc300)
	.awready (ds18_awready      ), // (axi_slave18) => (axi_monitor_s18,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds18_wid          ), // (axi_monitor_s18,axi_slave18) <= ()
	.wdata   (ds18_wdata        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wstrb   (ds18_wstrb        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wlast   (ds18_wlast        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wvalid  (ds18_wvalid       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wready  (ds18_wready       ), // (axi_slave18) => (axi_monitor_s18,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds18_bid          ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.bresp   (ds18_bresp        ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.bvalid  (ds18_bvalid       ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.bready  (ds18_bready       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds18_arid         ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.araddr  (ds18_araddr       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arlen   (ds18_arlen        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arsize  (ds18_arsize       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arburst (ds18_arburst      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arlock  ({1'b0,ds18_arlock}), // () <= ()
	.arcache (ds18_arcache      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arprot  (ds18_arprot       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arvalid (ds18_arvalid      ), // (axi_monitor_s18,axi_slave18,bench) <= (bmc300)
	.arready (ds18_arready      ), // (axi_slave18) => (axi_monitor_s18,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds18_rid          ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.rdata   (ds18_rdata        ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.rresp   (ds18_rresp        ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.rlast   (ds18_rlast        ), // (axi_slave18) => (axi_monitor_s18,bmc300)
	.rvalid  (ds18_rvalid       ), // (axi_slave18) => (axi_monitor_s18,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds18_rready       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave18) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave18

defparam axi_monitor_s18.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s18.AXI4 = 1'b1;
defparam axi_monitor_s18.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s18.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s18.MASTER_ID = 118;
defparam axi_monitor_s18.SLAVE_ID = 118;
axi_monitor axi_monitor_s18 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds18_awid         ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awaddr  (ds18_awaddr       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awlen   (ds18_awlen        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awsize  (ds18_awsize       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awburst (ds18_awburst      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awlock  ({1'b0,ds18_awlock}), // () <= ()
	.awcache (ds18_awcache      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awprot  (ds18_awprot       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.awvalid (ds18_awvalid      ), // (axi_monitor_s18,axi_slave18,bench) <= (bmc300)
	.awready (ds18_awready      ), // (axi_monitor_s18,bench,bmc300) <= (axi_slave18)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds18_wid          ), // (axi_monitor_s18,axi_slave18) <= ()
	.wdata   (ds18_wdata        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wstrb   (ds18_wstrb        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wlast   (ds18_wlast        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wvalid  (ds18_wvalid       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.wready  (ds18_wready       ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds18_bid          ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.bresp   (ds18_bresp        ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.bvalid  (ds18_bvalid       ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.bready  (ds18_bready       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds18_arid         ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.araddr  (ds18_araddr       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arlen   (ds18_arlen        ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arsize  (ds18_arsize       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arburst (ds18_arburst      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arlock  ({1'b0,ds18_arlock}), // () <= ()
	.arcache (ds18_arcache      ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arprot  (ds18_arprot       ), // (axi_monitor_s18,axi_slave18) <= (bmc300)
	.arvalid (ds18_arvalid      ), // (axi_monitor_s18,axi_slave18,bench) <= (bmc300)
	.arready (ds18_arready      ), // (axi_monitor_s18,bench,bmc300) <= (axi_slave18)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds18_rid          ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.rdata   (ds18_rdata        ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.rresp   (ds18_rresp        ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.rlast   (ds18_rlast        ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
	.rvalid  (ds18_rvalid       ), // (axi_monitor_s18,bmc300) <= (axi_slave18)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds18_rready       )  // (axi_monitor_s18,axi_slave18) <= (bmc300)
); // end of axi_monitor_s18

`endif // ATCBMC300_SLV18_SUPPORT
`ifdef ATCBMC300_SLV19_SUPPORT
defparam axi_slave19.ADDR_DECODE_WIDTH = `ATCBMC300_SLV19_SIZE+19;
defparam axi_slave19.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave19.AXI4 = 1'b1;
defparam axi_slave19.DATA_WIDTH = DATA_SIZE;
defparam axi_slave19.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave19.MEM_ADDR_WIDTH = `ATCBMC300_SLV19_SIZE+19;
defparam axi_slave19.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave19 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds19_awid         ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awaddr  (ds19_awaddr       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awlen   (ds19_awlen        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awsize  (ds19_awsize       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awburst (ds19_awburst      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awlock  ({1'b0,ds19_awlock}), // () <= ()
	.awcache (ds19_awcache      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awprot  (ds19_awprot       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awvalid (ds19_awvalid      ), // (axi_monitor_s19,axi_slave19,bench) <= (bmc300)
	.awready (ds19_awready      ), // (axi_slave19) => (axi_monitor_s19,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds19_wid          ), // (axi_monitor_s19,axi_slave19) <= ()
	.wdata   (ds19_wdata        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wstrb   (ds19_wstrb        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wlast   (ds19_wlast        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wvalid  (ds19_wvalid       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wready  (ds19_wready       ), // (axi_slave19) => (axi_monitor_s19,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds19_bid          ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.bresp   (ds19_bresp        ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.bvalid  (ds19_bvalid       ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.bready  (ds19_bready       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds19_arid         ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.araddr  (ds19_araddr       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arlen   (ds19_arlen        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arsize  (ds19_arsize       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arburst (ds19_arburst      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arlock  ({1'b0,ds19_arlock}), // () <= ()
	.arcache (ds19_arcache      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arprot  (ds19_arprot       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arvalid (ds19_arvalid      ), // (axi_monitor_s19,axi_slave19,bench) <= (bmc300)
	.arready (ds19_arready      ), // (axi_slave19) => (axi_monitor_s19,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds19_rid          ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.rdata   (ds19_rdata        ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.rresp   (ds19_rresp        ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.rlast   (ds19_rlast        ), // (axi_slave19) => (axi_monitor_s19,bmc300)
	.rvalid  (ds19_rvalid       ), // (axi_slave19) => (axi_monitor_s19,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds19_rready       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave19) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave19

defparam axi_monitor_s19.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s19.AXI4 = 1'b1;
defparam axi_monitor_s19.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s19.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s19.MASTER_ID = 119;
defparam axi_monitor_s19.SLAVE_ID = 119;
axi_monitor axi_monitor_s19 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds19_awid         ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awaddr  (ds19_awaddr       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awlen   (ds19_awlen        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awsize  (ds19_awsize       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awburst (ds19_awburst      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awlock  ({1'b0,ds19_awlock}), // () <= ()
	.awcache (ds19_awcache      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awprot  (ds19_awprot       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.awvalid (ds19_awvalid      ), // (axi_monitor_s19,axi_slave19,bench) <= (bmc300)
	.awready (ds19_awready      ), // (axi_monitor_s19,bench,bmc300) <= (axi_slave19)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds19_wid          ), // (axi_monitor_s19,axi_slave19) <= ()
	.wdata   (ds19_wdata        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wstrb   (ds19_wstrb        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wlast   (ds19_wlast        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wvalid  (ds19_wvalid       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.wready  (ds19_wready       ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds19_bid          ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.bresp   (ds19_bresp        ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.bvalid  (ds19_bvalid       ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.bready  (ds19_bready       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds19_arid         ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.araddr  (ds19_araddr       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arlen   (ds19_arlen        ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arsize  (ds19_arsize       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arburst (ds19_arburst      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arlock  ({1'b0,ds19_arlock}), // () <= ()
	.arcache (ds19_arcache      ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arprot  (ds19_arprot       ), // (axi_monitor_s19,axi_slave19) <= (bmc300)
	.arvalid (ds19_arvalid      ), // (axi_monitor_s19,axi_slave19,bench) <= (bmc300)
	.arready (ds19_arready      ), // (axi_monitor_s19,bench,bmc300) <= (axi_slave19)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds19_rid          ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.rdata   (ds19_rdata        ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.rresp   (ds19_rresp        ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.rlast   (ds19_rlast        ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
	.rvalid  (ds19_rvalid       ), // (axi_monitor_s19,bmc300) <= (axi_slave19)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds19_rready       )  // (axi_monitor_s19,axi_slave19) <= (bmc300)
); // end of axi_monitor_s19

`endif // ATCBMC300_SLV19_SUPPORT
`ifdef ATCBMC300_SLV20_SUPPORT
defparam axi_slave20.ADDR_DECODE_WIDTH = `ATCBMC300_SLV20_SIZE+19;
defparam axi_slave20.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave20.AXI4 = 1'b1;
defparam axi_slave20.DATA_WIDTH = DATA_SIZE;
defparam axi_slave20.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave20.MEM_ADDR_WIDTH = `ATCBMC300_SLV20_SIZE+19;
defparam axi_slave20.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave20 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds20_awid         ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awaddr  (ds20_awaddr       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awlen   (ds20_awlen        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awsize  (ds20_awsize       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awburst (ds20_awburst      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awlock  ({1'b0,ds20_awlock}), // () <= ()
	.awcache (ds20_awcache      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awprot  (ds20_awprot       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awvalid (ds20_awvalid      ), // (axi_monitor_s20,axi_slave20,bench) <= (bmc300)
	.awready (ds20_awready      ), // (axi_slave20) => (axi_monitor_s20,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds20_wid          ), // (axi_monitor_s20,axi_slave20) <= ()
	.wdata   (ds20_wdata        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wstrb   (ds20_wstrb        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wlast   (ds20_wlast        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wvalid  (ds20_wvalid       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wready  (ds20_wready       ), // (axi_slave20) => (axi_monitor_s20,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds20_bid          ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.bresp   (ds20_bresp        ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.bvalid  (ds20_bvalid       ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.bready  (ds20_bready       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds20_arid         ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.araddr  (ds20_araddr       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arlen   (ds20_arlen        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arsize  (ds20_arsize       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arburst (ds20_arburst      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arlock  ({1'b0,ds20_arlock}), // () <= ()
	.arcache (ds20_arcache      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arprot  (ds20_arprot       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arvalid (ds20_arvalid      ), // (axi_monitor_s20,axi_slave20,bench) <= (bmc300)
	.arready (ds20_arready      ), // (axi_slave20) => (axi_monitor_s20,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds20_rid          ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.rdata   (ds20_rdata        ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.rresp   (ds20_rresp        ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.rlast   (ds20_rlast        ), // (axi_slave20) => (axi_monitor_s20,bmc300)
	.rvalid  (ds20_rvalid       ), // (axi_slave20) => (axi_monitor_s20,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds20_rready       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave20) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave20

defparam axi_monitor_s20.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s20.AXI4 = 1'b1;
defparam axi_monitor_s20.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s20.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s20.MASTER_ID = 120;
defparam axi_monitor_s20.SLAVE_ID = 120;
axi_monitor axi_monitor_s20 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds20_awid         ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awaddr  (ds20_awaddr       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awlen   (ds20_awlen        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awsize  (ds20_awsize       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awburst (ds20_awburst      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awlock  ({1'b0,ds20_awlock}), // () <= ()
	.awcache (ds20_awcache      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awprot  (ds20_awprot       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.awvalid (ds20_awvalid      ), // (axi_monitor_s20,axi_slave20,bench) <= (bmc300)
	.awready (ds20_awready      ), // (axi_monitor_s20,bench,bmc300) <= (axi_slave20)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds20_wid          ), // (axi_monitor_s20,axi_slave20) <= ()
	.wdata   (ds20_wdata        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wstrb   (ds20_wstrb        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wlast   (ds20_wlast        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wvalid  (ds20_wvalid       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.wready  (ds20_wready       ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds20_bid          ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.bresp   (ds20_bresp        ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.bvalid  (ds20_bvalid       ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.bready  (ds20_bready       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds20_arid         ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.araddr  (ds20_araddr       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arlen   (ds20_arlen        ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arsize  (ds20_arsize       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arburst (ds20_arburst      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arlock  ({1'b0,ds20_arlock}), // () <= ()
	.arcache (ds20_arcache      ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arprot  (ds20_arprot       ), // (axi_monitor_s20,axi_slave20) <= (bmc300)
	.arvalid (ds20_arvalid      ), // (axi_monitor_s20,axi_slave20,bench) <= (bmc300)
	.arready (ds20_arready      ), // (axi_monitor_s20,bench,bmc300) <= (axi_slave20)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds20_rid          ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.rdata   (ds20_rdata        ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.rresp   (ds20_rresp        ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.rlast   (ds20_rlast        ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
	.rvalid  (ds20_rvalid       ), // (axi_monitor_s20,bmc300) <= (axi_slave20)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds20_rready       )  // (axi_monitor_s20,axi_slave20) <= (bmc300)
); // end of axi_monitor_s20

`endif // ATCBMC300_SLV20_SUPPORT
`ifdef ATCBMC300_SLV21_SUPPORT
defparam axi_slave21.ADDR_DECODE_WIDTH = `ATCBMC300_SLV21_SIZE+19;
defparam axi_slave21.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave21.AXI4 = 1'b1;
defparam axi_slave21.DATA_WIDTH = DATA_SIZE;
defparam axi_slave21.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave21.MEM_ADDR_WIDTH = `ATCBMC300_SLV21_SIZE+19;
defparam axi_slave21.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave21 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds21_awid         ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awaddr  (ds21_awaddr       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awlen   (ds21_awlen        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awsize  (ds21_awsize       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awburst (ds21_awburst      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awlock  ({1'b0,ds21_awlock}), // () <= ()
	.awcache (ds21_awcache      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awprot  (ds21_awprot       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awvalid (ds21_awvalid      ), // (axi_monitor_s21,axi_slave21,bench) <= (bmc300)
	.awready (ds21_awready      ), // (axi_slave21) => (axi_monitor_s21,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds21_wid          ), // (axi_monitor_s21,axi_slave21) <= ()
	.wdata   (ds21_wdata        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wstrb   (ds21_wstrb        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wlast   (ds21_wlast        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wvalid  (ds21_wvalid       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wready  (ds21_wready       ), // (axi_slave21) => (axi_monitor_s21,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds21_bid          ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.bresp   (ds21_bresp        ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.bvalid  (ds21_bvalid       ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.bready  (ds21_bready       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds21_arid         ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.araddr  (ds21_araddr       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arlen   (ds21_arlen        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arsize  (ds21_arsize       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arburst (ds21_arburst      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arlock  ({1'b0,ds21_arlock}), // () <= ()
	.arcache (ds21_arcache      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arprot  (ds21_arprot       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arvalid (ds21_arvalid      ), // (axi_monitor_s21,axi_slave21,bench) <= (bmc300)
	.arready (ds21_arready      ), // (axi_slave21) => (axi_monitor_s21,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds21_rid          ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.rdata   (ds21_rdata        ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.rresp   (ds21_rresp        ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.rlast   (ds21_rlast        ), // (axi_slave21) => (axi_monitor_s21,bmc300)
	.rvalid  (ds21_rvalid       ), // (axi_slave21) => (axi_monitor_s21,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds21_rready       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave21) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave21

defparam axi_monitor_s21.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s21.AXI4 = 1'b1;
defparam axi_monitor_s21.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s21.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s21.MASTER_ID = 121;
defparam axi_monitor_s21.SLAVE_ID = 121;
axi_monitor axi_monitor_s21 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds21_awid         ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awaddr  (ds21_awaddr       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awlen   (ds21_awlen        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awsize  (ds21_awsize       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awburst (ds21_awburst      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awlock  ({1'b0,ds21_awlock}), // () <= ()
	.awcache (ds21_awcache      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awprot  (ds21_awprot       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.awvalid (ds21_awvalid      ), // (axi_monitor_s21,axi_slave21,bench) <= (bmc300)
	.awready (ds21_awready      ), // (axi_monitor_s21,bench,bmc300) <= (axi_slave21)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds21_wid          ), // (axi_monitor_s21,axi_slave21) <= ()
	.wdata   (ds21_wdata        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wstrb   (ds21_wstrb        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wlast   (ds21_wlast        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wvalid  (ds21_wvalid       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.wready  (ds21_wready       ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds21_bid          ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.bresp   (ds21_bresp        ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.bvalid  (ds21_bvalid       ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.bready  (ds21_bready       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds21_arid         ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.araddr  (ds21_araddr       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arlen   (ds21_arlen        ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arsize  (ds21_arsize       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arburst (ds21_arburst      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arlock  ({1'b0,ds21_arlock}), // () <= ()
	.arcache (ds21_arcache      ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arprot  (ds21_arprot       ), // (axi_monitor_s21,axi_slave21) <= (bmc300)
	.arvalid (ds21_arvalid      ), // (axi_monitor_s21,axi_slave21,bench) <= (bmc300)
	.arready (ds21_arready      ), // (axi_monitor_s21,bench,bmc300) <= (axi_slave21)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds21_rid          ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.rdata   (ds21_rdata        ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.rresp   (ds21_rresp        ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.rlast   (ds21_rlast        ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
	.rvalid  (ds21_rvalid       ), // (axi_monitor_s21,bmc300) <= (axi_slave21)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds21_rready       )  // (axi_monitor_s21,axi_slave21) <= (bmc300)
); // end of axi_monitor_s21

`endif // ATCBMC300_SLV21_SUPPORT
`ifdef ATCBMC300_SLV22_SUPPORT
defparam axi_slave22.ADDR_DECODE_WIDTH = `ATCBMC300_SLV22_SIZE+19;
defparam axi_slave22.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave22.AXI4 = 1'b1;
defparam axi_slave22.DATA_WIDTH = DATA_SIZE;
defparam axi_slave22.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave22.MEM_ADDR_WIDTH = `ATCBMC300_SLV22_SIZE+19;
defparam axi_slave22.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave22 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds22_awid         ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awaddr  (ds22_awaddr       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awlen   (ds22_awlen        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awsize  (ds22_awsize       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awburst (ds22_awburst      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awlock  ({1'b0,ds22_awlock}), // () <= ()
	.awcache (ds22_awcache      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awprot  (ds22_awprot       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awvalid (ds22_awvalid      ), // (axi_monitor_s22,axi_slave22,bench) <= (bmc300)
	.awready (ds22_awready      ), // (axi_slave22) => (axi_monitor_s22,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds22_wid          ), // (axi_monitor_s22,axi_slave22) <= ()
	.wdata   (ds22_wdata        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wstrb   (ds22_wstrb        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wlast   (ds22_wlast        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wvalid  (ds22_wvalid       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wready  (ds22_wready       ), // (axi_slave22) => (axi_monitor_s22,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds22_bid          ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.bresp   (ds22_bresp        ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.bvalid  (ds22_bvalid       ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.bready  (ds22_bready       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds22_arid         ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.araddr  (ds22_araddr       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arlen   (ds22_arlen        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arsize  (ds22_arsize       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arburst (ds22_arburst      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arlock  ({1'b0,ds22_arlock}), // () <= ()
	.arcache (ds22_arcache      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arprot  (ds22_arprot       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arvalid (ds22_arvalid      ), // (axi_monitor_s22,axi_slave22,bench) <= (bmc300)
	.arready (ds22_arready      ), // (axi_slave22) => (axi_monitor_s22,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds22_rid          ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.rdata   (ds22_rdata        ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.rresp   (ds22_rresp        ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.rlast   (ds22_rlast        ), // (axi_slave22) => (axi_monitor_s22,bmc300)
	.rvalid  (ds22_rvalid       ), // (axi_slave22) => (axi_monitor_s22,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds22_rready       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave22) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave22

defparam axi_monitor_s22.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s22.AXI4 = 1'b1;
defparam axi_monitor_s22.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s22.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s22.MASTER_ID = 122;
defparam axi_monitor_s22.SLAVE_ID = 122;
axi_monitor axi_monitor_s22 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds22_awid         ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awaddr  (ds22_awaddr       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awlen   (ds22_awlen        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awsize  (ds22_awsize       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awburst (ds22_awburst      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awlock  ({1'b0,ds22_awlock}), // () <= ()
	.awcache (ds22_awcache      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awprot  (ds22_awprot       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.awvalid (ds22_awvalid      ), // (axi_monitor_s22,axi_slave22,bench) <= (bmc300)
	.awready (ds22_awready      ), // (axi_monitor_s22,bench,bmc300) <= (axi_slave22)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds22_wid          ), // (axi_monitor_s22,axi_slave22) <= ()
	.wdata   (ds22_wdata        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wstrb   (ds22_wstrb        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wlast   (ds22_wlast        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wvalid  (ds22_wvalid       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.wready  (ds22_wready       ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds22_bid          ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.bresp   (ds22_bresp        ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.bvalid  (ds22_bvalid       ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.bready  (ds22_bready       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds22_arid         ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.araddr  (ds22_araddr       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arlen   (ds22_arlen        ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arsize  (ds22_arsize       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arburst (ds22_arburst      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arlock  ({1'b0,ds22_arlock}), // () <= ()
	.arcache (ds22_arcache      ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arprot  (ds22_arprot       ), // (axi_monitor_s22,axi_slave22) <= (bmc300)
	.arvalid (ds22_arvalid      ), // (axi_monitor_s22,axi_slave22,bench) <= (bmc300)
	.arready (ds22_arready      ), // (axi_monitor_s22,bench,bmc300) <= (axi_slave22)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds22_rid          ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.rdata   (ds22_rdata        ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.rresp   (ds22_rresp        ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.rlast   (ds22_rlast        ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
	.rvalid  (ds22_rvalid       ), // (axi_monitor_s22,bmc300) <= (axi_slave22)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds22_rready       )  // (axi_monitor_s22,axi_slave22) <= (bmc300)
); // end of axi_monitor_s22

`endif // ATCBMC300_SLV22_SUPPORT
`ifdef ATCBMC300_SLV23_SUPPORT
defparam axi_slave23.ADDR_DECODE_WIDTH = `ATCBMC300_SLV23_SIZE+19;
defparam axi_slave23.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave23.AXI4 = 1'b1;
defparam axi_slave23.DATA_WIDTH = DATA_SIZE;
defparam axi_slave23.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave23.MEM_ADDR_WIDTH = `ATCBMC300_SLV23_SIZE+19;
defparam axi_slave23.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave23 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds23_awid         ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awaddr  (ds23_awaddr       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awlen   (ds23_awlen        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awsize  (ds23_awsize       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awburst (ds23_awburst      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awlock  ({1'b0,ds23_awlock}), // () <= ()
	.awcache (ds23_awcache      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awprot  (ds23_awprot       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awvalid (ds23_awvalid      ), // (axi_monitor_s23,axi_slave23,bench) <= (bmc300)
	.awready (ds23_awready      ), // (axi_slave23) => (axi_monitor_s23,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds23_wid          ), // (axi_monitor_s23,axi_slave23) <= ()
	.wdata   (ds23_wdata        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wstrb   (ds23_wstrb        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wlast   (ds23_wlast        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wvalid  (ds23_wvalid       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wready  (ds23_wready       ), // (axi_slave23) => (axi_monitor_s23,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds23_bid          ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.bresp   (ds23_bresp        ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.bvalid  (ds23_bvalid       ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.bready  (ds23_bready       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds23_arid         ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.araddr  (ds23_araddr       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arlen   (ds23_arlen        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arsize  (ds23_arsize       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arburst (ds23_arburst      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arlock  ({1'b0,ds23_arlock}), // () <= ()
	.arcache (ds23_arcache      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arprot  (ds23_arprot       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arvalid (ds23_arvalid      ), // (axi_monitor_s23,axi_slave23,bench) <= (bmc300)
	.arready (ds23_arready      ), // (axi_slave23) => (axi_monitor_s23,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds23_rid          ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.rdata   (ds23_rdata        ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.rresp   (ds23_rresp        ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.rlast   (ds23_rlast        ), // (axi_slave23) => (axi_monitor_s23,bmc300)
	.rvalid  (ds23_rvalid       ), // (axi_slave23) => (axi_monitor_s23,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds23_rready       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave23) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave23

defparam axi_monitor_s23.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s23.AXI4 = 1'b1;
defparam axi_monitor_s23.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s23.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s23.MASTER_ID = 123;
defparam axi_monitor_s23.SLAVE_ID = 123;
axi_monitor axi_monitor_s23 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds23_awid         ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awaddr  (ds23_awaddr       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awlen   (ds23_awlen        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awsize  (ds23_awsize       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awburst (ds23_awburst      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awlock  ({1'b0,ds23_awlock}), // () <= ()
	.awcache (ds23_awcache      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awprot  (ds23_awprot       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.awvalid (ds23_awvalid      ), // (axi_monitor_s23,axi_slave23,bench) <= (bmc300)
	.awready (ds23_awready      ), // (axi_monitor_s23,bench,bmc300) <= (axi_slave23)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds23_wid          ), // (axi_monitor_s23,axi_slave23) <= ()
	.wdata   (ds23_wdata        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wstrb   (ds23_wstrb        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wlast   (ds23_wlast        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wvalid  (ds23_wvalid       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.wready  (ds23_wready       ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds23_bid          ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.bresp   (ds23_bresp        ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.bvalid  (ds23_bvalid       ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.bready  (ds23_bready       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds23_arid         ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.araddr  (ds23_araddr       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arlen   (ds23_arlen        ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arsize  (ds23_arsize       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arburst (ds23_arburst      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arlock  ({1'b0,ds23_arlock}), // () <= ()
	.arcache (ds23_arcache      ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arprot  (ds23_arprot       ), // (axi_monitor_s23,axi_slave23) <= (bmc300)
	.arvalid (ds23_arvalid      ), // (axi_monitor_s23,axi_slave23,bench) <= (bmc300)
	.arready (ds23_arready      ), // (axi_monitor_s23,bench,bmc300) <= (axi_slave23)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds23_rid          ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.rdata   (ds23_rdata        ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.rresp   (ds23_rresp        ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.rlast   (ds23_rlast        ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
	.rvalid  (ds23_rvalid       ), // (axi_monitor_s23,bmc300) <= (axi_slave23)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds23_rready       )  // (axi_monitor_s23,axi_slave23) <= (bmc300)
); // end of axi_monitor_s23

`endif // ATCBMC300_SLV23_SUPPORT
`ifdef ATCBMC300_SLV24_SUPPORT
defparam axi_slave24.ADDR_DECODE_WIDTH = `ATCBMC300_SLV24_SIZE+19;
defparam axi_slave24.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave24.AXI4 = 1'b1;
defparam axi_slave24.DATA_WIDTH = DATA_SIZE;
defparam axi_slave24.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave24.MEM_ADDR_WIDTH = `ATCBMC300_SLV24_SIZE+19;
defparam axi_slave24.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave24 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds24_awid         ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awaddr  (ds24_awaddr       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awlen   (ds24_awlen        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awsize  (ds24_awsize       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awburst (ds24_awburst      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awlock  ({1'b0,ds24_awlock}), // () <= ()
	.awcache (ds24_awcache      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awprot  (ds24_awprot       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awvalid (ds24_awvalid      ), // (axi_monitor_s24,axi_slave24,bench) <= (bmc300)
	.awready (ds24_awready      ), // (axi_slave24) => (axi_monitor_s24,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds24_wid          ), // (axi_monitor_s24,axi_slave24) <= ()
	.wdata   (ds24_wdata        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wstrb   (ds24_wstrb        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wlast   (ds24_wlast        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wvalid  (ds24_wvalid       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wready  (ds24_wready       ), // (axi_slave24) => (axi_monitor_s24,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds24_bid          ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.bresp   (ds24_bresp        ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.bvalid  (ds24_bvalid       ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.bready  (ds24_bready       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds24_arid         ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.araddr  (ds24_araddr       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arlen   (ds24_arlen        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arsize  (ds24_arsize       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arburst (ds24_arburst      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arlock  ({1'b0,ds24_arlock}), // () <= ()
	.arcache (ds24_arcache      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arprot  (ds24_arprot       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arvalid (ds24_arvalid      ), // (axi_monitor_s24,axi_slave24,bench) <= (bmc300)
	.arready (ds24_arready      ), // (axi_slave24) => (axi_monitor_s24,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds24_rid          ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.rdata   (ds24_rdata        ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.rresp   (ds24_rresp        ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.rlast   (ds24_rlast        ), // (axi_slave24) => (axi_monitor_s24,bmc300)
	.rvalid  (ds24_rvalid       ), // (axi_slave24) => (axi_monitor_s24,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds24_rready       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave24) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave24

defparam axi_monitor_s24.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s24.AXI4 = 1'b1;
defparam axi_monitor_s24.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s24.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s24.MASTER_ID = 124;
defparam axi_monitor_s24.SLAVE_ID = 124;
axi_monitor axi_monitor_s24 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds24_awid         ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awaddr  (ds24_awaddr       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awlen   (ds24_awlen        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awsize  (ds24_awsize       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awburst (ds24_awburst      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awlock  ({1'b0,ds24_awlock}), // () <= ()
	.awcache (ds24_awcache      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awprot  (ds24_awprot       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.awvalid (ds24_awvalid      ), // (axi_monitor_s24,axi_slave24,bench) <= (bmc300)
	.awready (ds24_awready      ), // (axi_monitor_s24,bench,bmc300) <= (axi_slave24)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds24_wid          ), // (axi_monitor_s24,axi_slave24) <= ()
	.wdata   (ds24_wdata        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wstrb   (ds24_wstrb        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wlast   (ds24_wlast        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wvalid  (ds24_wvalid       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.wready  (ds24_wready       ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds24_bid          ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.bresp   (ds24_bresp        ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.bvalid  (ds24_bvalid       ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.bready  (ds24_bready       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds24_arid         ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.araddr  (ds24_araddr       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arlen   (ds24_arlen        ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arsize  (ds24_arsize       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arburst (ds24_arburst      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arlock  ({1'b0,ds24_arlock}), // () <= ()
	.arcache (ds24_arcache      ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arprot  (ds24_arprot       ), // (axi_monitor_s24,axi_slave24) <= (bmc300)
	.arvalid (ds24_arvalid      ), // (axi_monitor_s24,axi_slave24,bench) <= (bmc300)
	.arready (ds24_arready      ), // (axi_monitor_s24,bench,bmc300) <= (axi_slave24)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds24_rid          ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.rdata   (ds24_rdata        ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.rresp   (ds24_rresp        ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.rlast   (ds24_rlast        ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
	.rvalid  (ds24_rvalid       ), // (axi_monitor_s24,bmc300) <= (axi_slave24)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds24_rready       )  // (axi_monitor_s24,axi_slave24) <= (bmc300)
); // end of axi_monitor_s24

`endif // ATCBMC300_SLV24_SUPPORT
`ifdef ATCBMC300_SLV25_SUPPORT
defparam axi_slave25.ADDR_DECODE_WIDTH = `ATCBMC300_SLV25_SIZE+19;
defparam axi_slave25.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave25.AXI4 = 1'b1;
defparam axi_slave25.DATA_WIDTH = DATA_SIZE;
defparam axi_slave25.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave25.MEM_ADDR_WIDTH = `ATCBMC300_SLV25_SIZE+19;
defparam axi_slave25.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave25 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds25_awid         ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awaddr  (ds25_awaddr       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awlen   (ds25_awlen        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awsize  (ds25_awsize       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awburst (ds25_awburst      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awlock  ({1'b0,ds25_awlock}), // () <= ()
	.awcache (ds25_awcache      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awprot  (ds25_awprot       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awvalid (ds25_awvalid      ), // (axi_monitor_s25,axi_slave25,bench) <= (bmc300)
	.awready (ds25_awready      ), // (axi_slave25) => (axi_monitor_s25,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds25_wid          ), // (axi_monitor_s25,axi_slave25) <= ()
	.wdata   (ds25_wdata        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wstrb   (ds25_wstrb        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wlast   (ds25_wlast        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wvalid  (ds25_wvalid       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wready  (ds25_wready       ), // (axi_slave25) => (axi_monitor_s25,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds25_bid          ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.bresp   (ds25_bresp        ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.bvalid  (ds25_bvalid       ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.bready  (ds25_bready       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds25_arid         ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.araddr  (ds25_araddr       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arlen   (ds25_arlen        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arsize  (ds25_arsize       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arburst (ds25_arburst      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arlock  ({1'b0,ds25_arlock}), // () <= ()
	.arcache (ds25_arcache      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arprot  (ds25_arprot       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arvalid (ds25_arvalid      ), // (axi_monitor_s25,axi_slave25,bench) <= (bmc300)
	.arready (ds25_arready      ), // (axi_slave25) => (axi_monitor_s25,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds25_rid          ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.rdata   (ds25_rdata        ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.rresp   (ds25_rresp        ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.rlast   (ds25_rlast        ), // (axi_slave25) => (axi_monitor_s25,bmc300)
	.rvalid  (ds25_rvalid       ), // (axi_slave25) => (axi_monitor_s25,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds25_rready       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave25) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave25

defparam axi_monitor_s25.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s25.AXI4 = 1'b1;
defparam axi_monitor_s25.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s25.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s25.MASTER_ID = 125;
defparam axi_monitor_s25.SLAVE_ID = 125;
axi_monitor axi_monitor_s25 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds25_awid         ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awaddr  (ds25_awaddr       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awlen   (ds25_awlen        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awsize  (ds25_awsize       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awburst (ds25_awburst      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awlock  ({1'b0,ds25_awlock}), // () <= ()
	.awcache (ds25_awcache      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awprot  (ds25_awprot       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.awvalid (ds25_awvalid      ), // (axi_monitor_s25,axi_slave25,bench) <= (bmc300)
	.awready (ds25_awready      ), // (axi_monitor_s25,bench,bmc300) <= (axi_slave25)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds25_wid          ), // (axi_monitor_s25,axi_slave25) <= ()
	.wdata   (ds25_wdata        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wstrb   (ds25_wstrb        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wlast   (ds25_wlast        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wvalid  (ds25_wvalid       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.wready  (ds25_wready       ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds25_bid          ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.bresp   (ds25_bresp        ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.bvalid  (ds25_bvalid       ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.bready  (ds25_bready       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds25_arid         ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.araddr  (ds25_araddr       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arlen   (ds25_arlen        ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arsize  (ds25_arsize       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arburst (ds25_arburst      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arlock  ({1'b0,ds25_arlock}), // () <= ()
	.arcache (ds25_arcache      ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arprot  (ds25_arprot       ), // (axi_monitor_s25,axi_slave25) <= (bmc300)
	.arvalid (ds25_arvalid      ), // (axi_monitor_s25,axi_slave25,bench) <= (bmc300)
	.arready (ds25_arready      ), // (axi_monitor_s25,bench,bmc300) <= (axi_slave25)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds25_rid          ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.rdata   (ds25_rdata        ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.rresp   (ds25_rresp        ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.rlast   (ds25_rlast        ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
	.rvalid  (ds25_rvalid       ), // (axi_monitor_s25,bmc300) <= (axi_slave25)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds25_rready       )  // (axi_monitor_s25,axi_slave25) <= (bmc300)
); // end of axi_monitor_s25

`endif // ATCBMC300_SLV25_SUPPORT
`ifdef ATCBMC300_SLV26_SUPPORT
defparam axi_slave26.ADDR_DECODE_WIDTH = `ATCBMC300_SLV26_SIZE+19;
defparam axi_slave26.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave26.AXI4 = 1'b1;
defparam axi_slave26.DATA_WIDTH = DATA_SIZE;
defparam axi_slave26.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave26.MEM_ADDR_WIDTH = `ATCBMC300_SLV26_SIZE+19;
defparam axi_slave26.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave26 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds26_awid         ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awaddr  (ds26_awaddr       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awlen   (ds26_awlen        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awsize  (ds26_awsize       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awburst (ds26_awburst      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awlock  ({1'b0,ds26_awlock}), // () <= ()
	.awcache (ds26_awcache      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awprot  (ds26_awprot       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awvalid (ds26_awvalid      ), // (axi_monitor_s26,axi_slave26,bench) <= (bmc300)
	.awready (ds26_awready      ), // (axi_slave26) => (axi_monitor_s26,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds26_wid          ), // (axi_monitor_s26,axi_slave26) <= ()
	.wdata   (ds26_wdata        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wstrb   (ds26_wstrb        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wlast   (ds26_wlast        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wvalid  (ds26_wvalid       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wready  (ds26_wready       ), // (axi_slave26) => (axi_monitor_s26,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds26_bid          ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.bresp   (ds26_bresp        ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.bvalid  (ds26_bvalid       ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.bready  (ds26_bready       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds26_arid         ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.araddr  (ds26_araddr       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arlen   (ds26_arlen        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arsize  (ds26_arsize       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arburst (ds26_arburst      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arlock  ({1'b0,ds26_arlock}), // () <= ()
	.arcache (ds26_arcache      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arprot  (ds26_arprot       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arvalid (ds26_arvalid      ), // (axi_monitor_s26,axi_slave26,bench) <= (bmc300)
	.arready (ds26_arready      ), // (axi_slave26) => (axi_monitor_s26,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds26_rid          ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.rdata   (ds26_rdata        ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.rresp   (ds26_rresp        ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.rlast   (ds26_rlast        ), // (axi_slave26) => (axi_monitor_s26,bmc300)
	.rvalid  (ds26_rvalid       ), // (axi_slave26) => (axi_monitor_s26,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds26_rready       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave26) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave26

defparam axi_monitor_s26.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s26.AXI4 = 1'b1;
defparam axi_monitor_s26.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s26.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s26.MASTER_ID = 126;
defparam axi_monitor_s26.SLAVE_ID = 126;
axi_monitor axi_monitor_s26 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds26_awid         ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awaddr  (ds26_awaddr       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awlen   (ds26_awlen        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awsize  (ds26_awsize       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awburst (ds26_awburst      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awlock  ({1'b0,ds26_awlock}), // () <= ()
	.awcache (ds26_awcache      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awprot  (ds26_awprot       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.awvalid (ds26_awvalid      ), // (axi_monitor_s26,axi_slave26,bench) <= (bmc300)
	.awready (ds26_awready      ), // (axi_monitor_s26,bench,bmc300) <= (axi_slave26)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds26_wid          ), // (axi_monitor_s26,axi_slave26) <= ()
	.wdata   (ds26_wdata        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wstrb   (ds26_wstrb        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wlast   (ds26_wlast        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wvalid  (ds26_wvalid       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.wready  (ds26_wready       ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds26_bid          ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.bresp   (ds26_bresp        ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.bvalid  (ds26_bvalid       ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.bready  (ds26_bready       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds26_arid         ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.araddr  (ds26_araddr       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arlen   (ds26_arlen        ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arsize  (ds26_arsize       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arburst (ds26_arburst      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arlock  ({1'b0,ds26_arlock}), // () <= ()
	.arcache (ds26_arcache      ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arprot  (ds26_arprot       ), // (axi_monitor_s26,axi_slave26) <= (bmc300)
	.arvalid (ds26_arvalid      ), // (axi_monitor_s26,axi_slave26,bench) <= (bmc300)
	.arready (ds26_arready      ), // (axi_monitor_s26,bench,bmc300) <= (axi_slave26)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds26_rid          ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.rdata   (ds26_rdata        ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.rresp   (ds26_rresp        ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.rlast   (ds26_rlast        ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
	.rvalid  (ds26_rvalid       ), // (axi_monitor_s26,bmc300) <= (axi_slave26)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds26_rready       )  // (axi_monitor_s26,axi_slave26) <= (bmc300)
); // end of axi_monitor_s26

`endif // ATCBMC300_SLV26_SUPPORT
`ifdef ATCBMC300_SLV27_SUPPORT
defparam axi_slave27.ADDR_DECODE_WIDTH = `ATCBMC300_SLV27_SIZE+19;
defparam axi_slave27.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave27.AXI4 = 1'b1;
defparam axi_slave27.DATA_WIDTH = DATA_SIZE;
defparam axi_slave27.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave27.MEM_ADDR_WIDTH = `ATCBMC300_SLV27_SIZE+19;
defparam axi_slave27.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave27 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds27_awid         ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awaddr  (ds27_awaddr       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awlen   (ds27_awlen        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awsize  (ds27_awsize       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awburst (ds27_awburst      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awlock  ({1'b0,ds27_awlock}), // () <= ()
	.awcache (ds27_awcache      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awprot  (ds27_awprot       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awvalid (ds27_awvalid      ), // (axi_monitor_s27,axi_slave27,bench) <= (bmc300)
	.awready (ds27_awready      ), // (axi_slave27) => (axi_monitor_s27,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds27_wid          ), // (axi_monitor_s27,axi_slave27) <= ()
	.wdata   (ds27_wdata        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wstrb   (ds27_wstrb        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wlast   (ds27_wlast        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wvalid  (ds27_wvalid       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wready  (ds27_wready       ), // (axi_slave27) => (axi_monitor_s27,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds27_bid          ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.bresp   (ds27_bresp        ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.bvalid  (ds27_bvalid       ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.bready  (ds27_bready       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds27_arid         ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.araddr  (ds27_araddr       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arlen   (ds27_arlen        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arsize  (ds27_arsize       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arburst (ds27_arburst      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arlock  ({1'b0,ds27_arlock}), // () <= ()
	.arcache (ds27_arcache      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arprot  (ds27_arprot       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arvalid (ds27_arvalid      ), // (axi_monitor_s27,axi_slave27,bench) <= (bmc300)
	.arready (ds27_arready      ), // (axi_slave27) => (axi_monitor_s27,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds27_rid          ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.rdata   (ds27_rdata        ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.rresp   (ds27_rresp        ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.rlast   (ds27_rlast        ), // (axi_slave27) => (axi_monitor_s27,bmc300)
	.rvalid  (ds27_rvalid       ), // (axi_slave27) => (axi_monitor_s27,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds27_rready       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave27) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave27

defparam axi_monitor_s27.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s27.AXI4 = 1'b1;
defparam axi_monitor_s27.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s27.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s27.MASTER_ID = 127;
defparam axi_monitor_s27.SLAVE_ID = 127;
axi_monitor axi_monitor_s27 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds27_awid         ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awaddr  (ds27_awaddr       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awlen   (ds27_awlen        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awsize  (ds27_awsize       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awburst (ds27_awburst      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awlock  ({1'b0,ds27_awlock}), // () <= ()
	.awcache (ds27_awcache      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awprot  (ds27_awprot       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.awvalid (ds27_awvalid      ), // (axi_monitor_s27,axi_slave27,bench) <= (bmc300)
	.awready (ds27_awready      ), // (axi_monitor_s27,bench,bmc300) <= (axi_slave27)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds27_wid          ), // (axi_monitor_s27,axi_slave27) <= ()
	.wdata   (ds27_wdata        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wstrb   (ds27_wstrb        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wlast   (ds27_wlast        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wvalid  (ds27_wvalid       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.wready  (ds27_wready       ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds27_bid          ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.bresp   (ds27_bresp        ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.bvalid  (ds27_bvalid       ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.bready  (ds27_bready       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds27_arid         ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.araddr  (ds27_araddr       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arlen   (ds27_arlen        ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arsize  (ds27_arsize       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arburst (ds27_arburst      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arlock  ({1'b0,ds27_arlock}), // () <= ()
	.arcache (ds27_arcache      ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arprot  (ds27_arprot       ), // (axi_monitor_s27,axi_slave27) <= (bmc300)
	.arvalid (ds27_arvalid      ), // (axi_monitor_s27,axi_slave27,bench) <= (bmc300)
	.arready (ds27_arready      ), // (axi_monitor_s27,bench,bmc300) <= (axi_slave27)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds27_rid          ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.rdata   (ds27_rdata        ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.rresp   (ds27_rresp        ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.rlast   (ds27_rlast        ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
	.rvalid  (ds27_rvalid       ), // (axi_monitor_s27,bmc300) <= (axi_slave27)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds27_rready       )  // (axi_monitor_s27,axi_slave27) <= (bmc300)
); // end of axi_monitor_s27

`endif // ATCBMC300_SLV27_SUPPORT
`ifdef ATCBMC300_SLV28_SUPPORT
defparam axi_slave28.ADDR_DECODE_WIDTH = `ATCBMC300_SLV28_SIZE+19;
defparam axi_slave28.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave28.AXI4 = 1'b1;
defparam axi_slave28.DATA_WIDTH = DATA_SIZE;
defparam axi_slave28.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave28.MEM_ADDR_WIDTH = `ATCBMC300_SLV28_SIZE+19;
defparam axi_slave28.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave28 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds28_awid         ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awaddr  (ds28_awaddr       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awlen   (ds28_awlen        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awsize  (ds28_awsize       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awburst (ds28_awburst      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awlock  ({1'b0,ds28_awlock}), // () <= ()
	.awcache (ds28_awcache      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awprot  (ds28_awprot       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awvalid (ds28_awvalid      ), // (axi_monitor_s28,axi_slave28,bench) <= (bmc300)
	.awready (ds28_awready      ), // (axi_slave28) => (axi_monitor_s28,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds28_wid          ), // (axi_monitor_s28,axi_slave28) <= ()
	.wdata   (ds28_wdata        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wstrb   (ds28_wstrb        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wlast   (ds28_wlast        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wvalid  (ds28_wvalid       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wready  (ds28_wready       ), // (axi_slave28) => (axi_monitor_s28,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds28_bid          ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.bresp   (ds28_bresp        ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.bvalid  (ds28_bvalid       ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.bready  (ds28_bready       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds28_arid         ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.araddr  (ds28_araddr       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arlen   (ds28_arlen        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arsize  (ds28_arsize       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arburst (ds28_arburst      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arlock  ({1'b0,ds28_arlock}), // () <= ()
	.arcache (ds28_arcache      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arprot  (ds28_arprot       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arvalid (ds28_arvalid      ), // (axi_monitor_s28,axi_slave28,bench) <= (bmc300)
	.arready (ds28_arready      ), // (axi_slave28) => (axi_monitor_s28,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds28_rid          ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.rdata   (ds28_rdata        ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.rresp   (ds28_rresp        ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.rlast   (ds28_rlast        ), // (axi_slave28) => (axi_monitor_s28,bmc300)
	.rvalid  (ds28_rvalid       ), // (axi_slave28) => (axi_monitor_s28,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds28_rready       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave28) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave28

defparam axi_monitor_s28.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s28.AXI4 = 1'b1;
defparam axi_monitor_s28.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s28.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s28.MASTER_ID = 128;
defparam axi_monitor_s28.SLAVE_ID = 128;
axi_monitor axi_monitor_s28 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds28_awid         ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awaddr  (ds28_awaddr       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awlen   (ds28_awlen        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awsize  (ds28_awsize       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awburst (ds28_awburst      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awlock  ({1'b0,ds28_awlock}), // () <= ()
	.awcache (ds28_awcache      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awprot  (ds28_awprot       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.awvalid (ds28_awvalid      ), // (axi_monitor_s28,axi_slave28,bench) <= (bmc300)
	.awready (ds28_awready      ), // (axi_monitor_s28,bench,bmc300) <= (axi_slave28)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds28_wid          ), // (axi_monitor_s28,axi_slave28) <= ()
	.wdata   (ds28_wdata        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wstrb   (ds28_wstrb        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wlast   (ds28_wlast        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wvalid  (ds28_wvalid       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.wready  (ds28_wready       ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds28_bid          ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.bresp   (ds28_bresp        ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.bvalid  (ds28_bvalid       ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.bready  (ds28_bready       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds28_arid         ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.araddr  (ds28_araddr       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arlen   (ds28_arlen        ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arsize  (ds28_arsize       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arburst (ds28_arburst      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arlock  ({1'b0,ds28_arlock}), // () <= ()
	.arcache (ds28_arcache      ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arprot  (ds28_arprot       ), // (axi_monitor_s28,axi_slave28) <= (bmc300)
	.arvalid (ds28_arvalid      ), // (axi_monitor_s28,axi_slave28,bench) <= (bmc300)
	.arready (ds28_arready      ), // (axi_monitor_s28,bench,bmc300) <= (axi_slave28)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds28_rid          ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.rdata   (ds28_rdata        ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.rresp   (ds28_rresp        ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.rlast   (ds28_rlast        ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
	.rvalid  (ds28_rvalid       ), // (axi_monitor_s28,bmc300) <= (axi_slave28)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds28_rready       )  // (axi_monitor_s28,axi_slave28) <= (bmc300)
); // end of axi_monitor_s28

`endif // ATCBMC300_SLV28_SUPPORT
`ifdef ATCBMC300_SLV29_SUPPORT
defparam axi_slave29.ADDR_DECODE_WIDTH = `ATCBMC300_SLV29_SIZE+19;
defparam axi_slave29.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave29.AXI4 = 1'b1;
defparam axi_slave29.DATA_WIDTH = DATA_SIZE;
defparam axi_slave29.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave29.MEM_ADDR_WIDTH = `ATCBMC300_SLV29_SIZE+19;
defparam axi_slave29.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave29 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds29_awid         ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awaddr  (ds29_awaddr       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awlen   (ds29_awlen        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awsize  (ds29_awsize       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awburst (ds29_awburst      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awlock  ({1'b0,ds29_awlock}), // () <= ()
	.awcache (ds29_awcache      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awprot  (ds29_awprot       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awvalid (ds29_awvalid      ), // (axi_monitor_s29,axi_slave29,bench) <= (bmc300)
	.awready (ds29_awready      ), // (axi_slave29) => (axi_monitor_s29,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds29_wid          ), // (axi_monitor_s29,axi_slave29) <= ()
	.wdata   (ds29_wdata        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wstrb   (ds29_wstrb        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wlast   (ds29_wlast        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wvalid  (ds29_wvalid       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wready  (ds29_wready       ), // (axi_slave29) => (axi_monitor_s29,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds29_bid          ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.bresp   (ds29_bresp        ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.bvalid  (ds29_bvalid       ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.bready  (ds29_bready       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds29_arid         ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.araddr  (ds29_araddr       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arlen   (ds29_arlen        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arsize  (ds29_arsize       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arburst (ds29_arburst      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arlock  ({1'b0,ds29_arlock}), // () <= ()
	.arcache (ds29_arcache      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arprot  (ds29_arprot       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arvalid (ds29_arvalid      ), // (axi_monitor_s29,axi_slave29,bench) <= (bmc300)
	.arready (ds29_arready      ), // (axi_slave29) => (axi_monitor_s29,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds29_rid          ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.rdata   (ds29_rdata        ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.rresp   (ds29_rresp        ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.rlast   (ds29_rlast        ), // (axi_slave29) => (axi_monitor_s29,bmc300)
	.rvalid  (ds29_rvalid       ), // (axi_slave29) => (axi_monitor_s29,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds29_rready       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave29) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave29

defparam axi_monitor_s29.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s29.AXI4 = 1'b1;
defparam axi_monitor_s29.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s29.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s29.MASTER_ID = 129;
defparam axi_monitor_s29.SLAVE_ID = 129;
axi_monitor axi_monitor_s29 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds29_awid         ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awaddr  (ds29_awaddr       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awlen   (ds29_awlen        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awsize  (ds29_awsize       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awburst (ds29_awburst      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awlock  ({1'b0,ds29_awlock}), // () <= ()
	.awcache (ds29_awcache      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awprot  (ds29_awprot       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.awvalid (ds29_awvalid      ), // (axi_monitor_s29,axi_slave29,bench) <= (bmc300)
	.awready (ds29_awready      ), // (axi_monitor_s29,bench,bmc300) <= (axi_slave29)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds29_wid          ), // (axi_monitor_s29,axi_slave29) <= ()
	.wdata   (ds29_wdata        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wstrb   (ds29_wstrb        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wlast   (ds29_wlast        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wvalid  (ds29_wvalid       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.wready  (ds29_wready       ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds29_bid          ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.bresp   (ds29_bresp        ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.bvalid  (ds29_bvalid       ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.bready  (ds29_bready       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds29_arid         ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.araddr  (ds29_araddr       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arlen   (ds29_arlen        ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arsize  (ds29_arsize       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arburst (ds29_arburst      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arlock  ({1'b0,ds29_arlock}), // () <= ()
	.arcache (ds29_arcache      ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arprot  (ds29_arprot       ), // (axi_monitor_s29,axi_slave29) <= (bmc300)
	.arvalid (ds29_arvalid      ), // (axi_monitor_s29,axi_slave29,bench) <= (bmc300)
	.arready (ds29_arready      ), // (axi_monitor_s29,bench,bmc300) <= (axi_slave29)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds29_rid          ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.rdata   (ds29_rdata        ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.rresp   (ds29_rresp        ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.rlast   (ds29_rlast        ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
	.rvalid  (ds29_rvalid       ), // (axi_monitor_s29,bmc300) <= (axi_slave29)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds29_rready       )  // (axi_monitor_s29,axi_slave29) <= (bmc300)
); // end of axi_monitor_s29

`endif // ATCBMC300_SLV29_SUPPORT
`ifdef ATCBMC300_SLV30_SUPPORT
defparam axi_slave30.ADDR_DECODE_WIDTH = `ATCBMC300_SLV30_SIZE+19;
defparam axi_slave30.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave30.AXI4 = 1'b1;
defparam axi_slave30.DATA_WIDTH = DATA_SIZE;
defparam axi_slave30.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave30.MEM_ADDR_WIDTH = `ATCBMC300_SLV30_SIZE+19;
defparam axi_slave30.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave30 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds30_awid         ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awaddr  (ds30_awaddr       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awlen   (ds30_awlen        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awsize  (ds30_awsize       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awburst (ds30_awburst      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awlock  ({1'b0,ds30_awlock}), // () <= ()
	.awcache (ds30_awcache      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awprot  (ds30_awprot       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awvalid (ds30_awvalid      ), // (axi_monitor_s30,axi_slave30,bench) <= (bmc300)
	.awready (ds30_awready      ), // (axi_slave30) => (axi_monitor_s30,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds30_wid          ), // (axi_monitor_s30,axi_slave30) <= ()
	.wdata   (ds30_wdata        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wstrb   (ds30_wstrb        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wlast   (ds30_wlast        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wvalid  (ds30_wvalid       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wready  (ds30_wready       ), // (axi_slave30) => (axi_monitor_s30,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds30_bid          ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.bresp   (ds30_bresp        ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.bvalid  (ds30_bvalid       ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.bready  (ds30_bready       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds30_arid         ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.araddr  (ds30_araddr       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arlen   (ds30_arlen        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arsize  (ds30_arsize       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arburst (ds30_arburst      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arlock  ({1'b0,ds30_arlock}), // () <= ()
	.arcache (ds30_arcache      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arprot  (ds30_arprot       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arvalid (ds30_arvalid      ), // (axi_monitor_s30,axi_slave30,bench) <= (bmc300)
	.arready (ds30_arready      ), // (axi_slave30) => (axi_monitor_s30,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds30_rid          ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.rdata   (ds30_rdata        ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.rresp   (ds30_rresp        ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.rlast   (ds30_rlast        ), // (axi_slave30) => (axi_monitor_s30,bmc300)
	.rvalid  (ds30_rvalid       ), // (axi_slave30) => (axi_monitor_s30,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds30_rready       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave30) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave30

defparam axi_monitor_s30.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s30.AXI4 = 1'b1;
defparam axi_monitor_s30.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s30.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s30.MASTER_ID = 130;
defparam axi_monitor_s30.SLAVE_ID = 130;
axi_monitor axi_monitor_s30 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds30_awid         ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awaddr  (ds30_awaddr       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awlen   (ds30_awlen        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awsize  (ds30_awsize       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awburst (ds30_awburst      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awlock  ({1'b0,ds30_awlock}), // () <= ()
	.awcache (ds30_awcache      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awprot  (ds30_awprot       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.awvalid (ds30_awvalid      ), // (axi_monitor_s30,axi_slave30,bench) <= (bmc300)
	.awready (ds30_awready      ), // (axi_monitor_s30,bench,bmc300) <= (axi_slave30)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds30_wid          ), // (axi_monitor_s30,axi_slave30) <= ()
	.wdata   (ds30_wdata        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wstrb   (ds30_wstrb        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wlast   (ds30_wlast        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wvalid  (ds30_wvalid       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.wready  (ds30_wready       ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds30_bid          ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.bresp   (ds30_bresp        ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.bvalid  (ds30_bvalid       ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.bready  (ds30_bready       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds30_arid         ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.araddr  (ds30_araddr       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arlen   (ds30_arlen        ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arsize  (ds30_arsize       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arburst (ds30_arburst      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arlock  ({1'b0,ds30_arlock}), // () <= ()
	.arcache (ds30_arcache      ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arprot  (ds30_arprot       ), // (axi_monitor_s30,axi_slave30) <= (bmc300)
	.arvalid (ds30_arvalid      ), // (axi_monitor_s30,axi_slave30,bench) <= (bmc300)
	.arready (ds30_arready      ), // (axi_monitor_s30,bench,bmc300) <= (axi_slave30)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds30_rid          ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.rdata   (ds30_rdata        ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.rresp   (ds30_rresp        ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.rlast   (ds30_rlast        ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
	.rvalid  (ds30_rvalid       ), // (axi_monitor_s30,bmc300) <= (axi_slave30)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds30_rready       )  // (axi_monitor_s30,axi_slave30) <= (bmc300)
); // end of axi_monitor_s30

`endif // ATCBMC300_SLV30_SUPPORT
`ifdef ATCBMC300_SLV31_SUPPORT
defparam axi_slave31.ADDR_DECODE_WIDTH = `ATCBMC300_SLV31_SIZE+19;
defparam axi_slave31.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_slave31.AXI4 = 1'b1;
defparam axi_slave31.DATA_WIDTH = DATA_SIZE;
defparam axi_slave31.ID_WIDTH = DS_ID_WIDTH;
defparam axi_slave31.MEM_ADDR_WIDTH = `ATCBMC300_SLV31_SIZE+19;
defparam axi_slave31.RAND_INIT_ON_READ_X = 1'b1;
axi_slave_model axi_slave31 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds31_awid         ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awaddr  (ds31_awaddr       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awlen   (ds31_awlen        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awsize  (ds31_awsize       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awburst (ds31_awburst      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awlock  ({1'b0,ds31_awlock}), // () <= ()
	.awcache (ds31_awcache      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awprot  (ds31_awprot       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awvalid (ds31_awvalid      ), // (axi_monitor_s31,axi_slave31,bench) <= (bmc300)
	.awready (ds31_awready      ), // (axi_slave31) => (axi_monitor_s31,bench,bmc300)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds31_wid          ), // (axi_monitor_s31,axi_slave31) <= ()
	.wdata   (ds31_wdata        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wstrb   (ds31_wstrb        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wlast   (ds31_wlast        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wvalid  (ds31_wvalid       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wready  (ds31_wready       ), // (axi_slave31) => (axi_monitor_s31,bmc300)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds31_bid          ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.bresp   (ds31_bresp        ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.bvalid  (ds31_bvalid       ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.bready  (ds31_bready       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds31_arid         ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.araddr  (ds31_araddr       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arlen   (ds31_arlen        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arsize  (ds31_arsize       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arburst (ds31_arburst      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arlock  ({1'b0,ds31_arlock}), // () <= ()
	.arcache (ds31_arcache      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arprot  (ds31_arprot       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arvalid (ds31_arvalid      ), // (axi_monitor_s31,axi_slave31,bench) <= (bmc300)
	.arready (ds31_arready      ), // (axi_slave31) => (axi_monitor_s31,bench,bmc300)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds31_rid          ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.rdata   (ds31_rdata        ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.rresp   (ds31_rresp        ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.rlast   (ds31_rlast        ), // (axi_slave31) => (axi_monitor_s31,bmc300)
	.rvalid  (ds31_rvalid       ), // (axi_slave31) => (axi_monitor_s31,bmc300)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds31_rready       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.csysreq (1'b0              ), // (axi_slave31) <= ()
	.csysack (                  ), // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
	.cactive (                  )  // (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) => ()
); // end of axi_slave31

defparam axi_monitor_s31.ADDR_WIDTH = ADDR_WIDTH;
defparam axi_monitor_s31.AXI4 = 1'b1;
defparam axi_monitor_s31.DATA_WIDTH = DATA_SIZE;
defparam axi_monitor_s31.ID_WIDTH = DS_ID_WIDTH;
defparam axi_monitor_s31.MASTER_ID = 131;
defparam axi_monitor_s31.SLAVE_ID = 131;
axi_monitor axi_monitor_s31 (
	.aclk    (aclk              ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.aresetn (aresetn           ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9,bmc300) <= (bench)
	.awid    (ds31_awid         ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awaddr  (ds31_awaddr       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awlen   (ds31_awlen        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awsize  (ds31_awsize       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awburst (ds31_awburst      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awlock  ({1'b0,ds31_awlock}), // () <= ()
	.awcache (ds31_awcache      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awprot  (ds31_awprot       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.awvalid (ds31_awvalid      ), // (axi_monitor_s31,axi_slave31,bench) <= (bmc300)
	.awready (ds31_awready      ), // (axi_monitor_s31,bench,bmc300) <= (axi_slave31)
   `ifdef NDS_AXI_AWREGION_SUPPORT
	.awregion(awregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWREGION_SUPPORT
   `ifdef NDS_AXI_AWQOS_SUPPORT
	.awqos   (awqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWQOS_SUPPORT
   `ifdef NDS_AXI_AWUSER_SUPPORT
	.awuser  (awuser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_AWUSER_SUPPORT
	.wid     (ds31_wid          ), // (axi_monitor_s31,axi_slave31) <= ()
	.wdata   (ds31_wdata        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wstrb   (ds31_wstrb        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wlast   (ds31_wlast        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wvalid  (ds31_wvalid       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.wready  (ds31_wready       ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
   `ifdef NDS_AXI_WUSER_SUPPORT
	.wuser   (wuser             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_WUSER_SUPPORT
	.bid     (ds31_bid          ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.bresp   (ds31_bresp        ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.bvalid  (ds31_bvalid       ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.bready  (ds31_bready       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
   `ifdef NDS_AXI_BUSER_SUPPORT
	.buser   (buser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_BUSER_SUPPORT
	.arid    (ds31_arid         ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.araddr  (ds31_araddr       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arlen   (ds31_arlen        ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arsize  (ds31_arsize       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arburst (ds31_arburst      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arlock  ({1'b0,ds31_arlock}), // () <= ()
	.arcache (ds31_arcache      ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arprot  (ds31_arprot       ), // (axi_monitor_s31,axi_slave31) <= (bmc300)
	.arvalid (ds31_arvalid      ), // (axi_monitor_s31,axi_slave31,bench) <= (bmc300)
	.arready (ds31_arready      ), // (axi_monitor_s31,bench,bmc300) <= (axi_slave31)
   `ifdef NDS_AXI_ARREGION_SUPPORT
	.arregion(arregion          ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARREGION_SUPPORT
   `ifdef NDS_AXI_ARQOS_SUPPORT
	.arqos   (arqos             ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARQOS_SUPPORT
   `ifdef NDS_AXI_ARUSER_SUPPORT
	.aruser  (aruser            ), // (axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9,axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9) <= (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9)
   `endif // NDS_AXI_ARUSER_SUPPORT
	.rid     (ds31_rid          ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.rdata   (ds31_rdata        ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.rresp   (ds31_rresp        ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.rlast   (ds31_rlast        ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
	.rvalid  (ds31_rvalid       ), // (axi_monitor_s31,bmc300) <= (axi_slave31)
   `ifdef NDS_AXI_RUSER_SUPPORT
	.ruser   (ruser             ), // (axi_master0,axi_master1,axi_master10,axi_master11,axi_master12,axi_master13,axi_master14,axi_master15,axi_master2,axi_master3,axi_master4,axi_master5,axi_master6,axi_master7,axi_master8,axi_master9,axi_monitor_m0,axi_monitor_m1,axi_monitor_m10,axi_monitor_m11,axi_monitor_m12,axi_monitor_m13,axi_monitor_m14,axi_monitor_m15,axi_monitor_m2,axi_monitor_m3,axi_monitor_m4,axi_monitor_m5,axi_monitor_m6,axi_monitor_m7,axi_monitor_m8,axi_monitor_m9,axi_monitor_s1,axi_monitor_s10,axi_monitor_s11,axi_monitor_s12,axi_monitor_s13,axi_monitor_s14,axi_monitor_s15,axi_monitor_s16,axi_monitor_s17,axi_monitor_s18,axi_monitor_s19,axi_monitor_s2,axi_monitor_s20,axi_monitor_s21,axi_monitor_s22,axi_monitor_s23,axi_monitor_s24,axi_monitor_s25,axi_monitor_s26,axi_monitor_s27,axi_monitor_s28,axi_monitor_s29,axi_monitor_s3,axi_monitor_s30,axi_monitor_s31,axi_monitor_s4,axi_monitor_s5,axi_monitor_s6,axi_monitor_s7,axi_monitor_s8,axi_monitor_s9) <= (axi_slave1,axi_slave10,axi_slave11,axi_slave12,axi_slave13,axi_slave14,axi_slave15,axi_slave16,axi_slave17,axi_slave18,axi_slave19,axi_slave2,axi_slave20,axi_slave21,axi_slave22,axi_slave23,axi_slave24,axi_slave25,axi_slave26,axi_slave27,axi_slave28,axi_slave29,axi_slave3,axi_slave30,axi_slave31,axi_slave4,axi_slave5,axi_slave6,axi_slave7,axi_slave8,axi_slave9)
   `endif // NDS_AXI_RUSER_SUPPORT
	.rready  (ds31_rready       )  // (axi_monitor_s31,axi_slave31) <= (bmc300)
); // end of axi_monitor_s31

`endif // ATCBMC300_SLV31_SUPPORT
endmodule
`ifdef NDS_SCOREBOARD_EN
`ifdef ATCBMC300_MST0_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master0 scb_axim_mon scb_axim_mon (.*, .model_id(8'd0));
`endif
`ifdef ATCBMC300_MST1_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master1 scb_axim_mon scb_axim_mon (.*, .model_id(8'd1));
`endif
`ifdef ATCBMC300_MST2_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master2 scb_axim_mon scb_axim_mon (.*, .model_id(8'd2));
`endif
`ifdef ATCBMC300_MST3_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master3 scb_axim_mon scb_axim_mon (.*, .model_id(8'd3));
`endif
`ifdef ATCBMC300_MST4_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master4 scb_axim_mon scb_axim_mon (.*, .model_id(8'd4));
`endif
`ifdef ATCBMC300_MST5_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master5 scb_axim_mon scb_axim_mon (.*, .model_id(8'd5));
`endif
`ifdef ATCBMC300_MST6_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master6 scb_axim_mon scb_axim_mon (.*, .model_id(8'd6));
`endif
`ifdef ATCBMC300_MST7_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master7 scb_axim_mon scb_axim_mon (.*, .model_id(8'd7));
`endif
`ifdef ATCBMC300_MST8_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master8 scb_axim_mon scb_axim_mon (.*, .model_id(8'd8));
`endif
`ifdef ATCBMC300_MST9_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master9 scb_axim_mon scb_axim_mon (.*, .model_id(8'd9));
`endif
`ifdef ATCBMC300_MST10_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master10 scb_axim_mon scb_axim_mon (.*, .model_id(8'd10));
`endif
`ifdef ATCBMC300_MST11_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master11 scb_axim_mon scb_axim_mon (.*, .model_id(8'd11));
`endif
`ifdef ATCBMC300_MST12_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master12 scb_axim_mon scb_axim_mon (.*, .model_id(8'd12));
`endif
`ifdef ATCBMC300_MST13_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master13 scb_axim_mon scb_axim_mon (.*, .model_id(8'd13));
`endif
`ifdef ATCBMC300_MST14_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master14 scb_axim_mon scb_axim_mon (.*, .model_id(8'd14));
`endif
`ifdef ATCBMC300_MST15_SUPPORT
bind axi_master_model :`NDS_SYSTEM.axi_master15 scb_axim_mon scb_axim_mon (.*, .model_id(8'd15));
`endif

`ifdef ATCBMC300_SLV1_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave1 scb_axis_mon scb_axis_mon (.*, .model_id(8'd1));
`endif
`ifdef ATCBMC300_SLV2_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave2 scb_axis_mon scb_axis_mon (.*, .model_id(8'd2));
`endif
`ifdef ATCBMC300_SLV3_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave3 scb_axis_mon scb_axis_mon (.*, .model_id(8'd3));
`endif
`ifdef ATCBMC300_SLV4_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave4 scb_axis_mon scb_axis_mon (.*, .model_id(8'd4));
`endif
`ifdef ATCBMC300_SLV5_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave5 scb_axis_mon scb_axis_mon (.*, .model_id(8'd5));
`endif
`ifdef ATCBMC300_SLV6_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave6 scb_axis_mon scb_axis_mon (.*, .model_id(8'd6));
`endif
`ifdef ATCBMC300_SLV7_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave7 scb_axis_mon scb_axis_mon (.*, .model_id(8'd7));
`endif
`ifdef ATCBMC300_SLV8_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave8 scb_axis_mon scb_axis_mon (.*, .model_id(8'd8));
`endif
`ifdef ATCBMC300_SLV9_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave9 scb_axis_mon scb_axis_mon (.*, .model_id(8'd9));
`endif
`ifdef ATCBMC300_SLV10_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave10 scb_axis_mon scb_axis_mon (.*, .model_id(8'd10));
`endif
`ifdef ATCBMC300_SLV11_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave11 scb_axis_mon scb_axis_mon (.*, .model_id(8'd11));
`endif
`ifdef ATCBMC300_SLV12_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave12 scb_axis_mon scb_axis_mon (.*, .model_id(8'd12));
`endif
`ifdef ATCBMC300_SLV13_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave13 scb_axis_mon scb_axis_mon (.*, .model_id(8'd13));
`endif
`ifdef ATCBMC300_SLV14_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave14 scb_axis_mon scb_axis_mon (.*, .model_id(8'd14));
`endif
`ifdef ATCBMC300_SLV15_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave15 scb_axis_mon scb_axis_mon (.*, .model_id(8'd15));
`endif
`ifdef ATCBMC300_SLV16_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave16 scb_axis_mon scb_axis_mon (.*, .model_id(8'd16));
`endif
`ifdef ATCBMC300_SLV17_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave17 scb_axis_mon scb_axis_mon (.*, .model_id(8'd17));
`endif
`ifdef ATCBMC300_SLV18_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave18 scb_axis_mon scb_axis_mon (.*, .model_id(8'd18));
`endif
`ifdef ATCBMC300_SLV19_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave19 scb_axis_mon scb_axis_mon (.*, .model_id(8'd19));
`endif
`ifdef ATCBMC300_SLV20_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave20 scb_axis_mon scb_axis_mon (.*, .model_id(8'd20));
`endif
`ifdef ATCBMC300_SLV21_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave21 scb_axis_mon scb_axis_mon (.*, .model_id(8'd21));
`endif
`ifdef ATCBMC300_SLV22_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave22 scb_axis_mon scb_axis_mon (.*, .model_id(8'd22));
`endif
`ifdef ATCBMC300_SLV23_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave23 scb_axis_mon scb_axis_mon (.*, .model_id(8'd23));
`endif
`ifdef ATCBMC300_SLV24_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave24 scb_axis_mon scb_axis_mon (.*, .model_id(8'd24));
`endif
`ifdef ATCBMC300_SLV25_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave25 scb_axis_mon scb_axis_mon (.*, .model_id(8'd25));
`endif
`ifdef ATCBMC300_SLV26_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave26 scb_axis_mon scb_axis_mon (.*, .model_id(8'd26));
`endif
`ifdef ATCBMC300_SLV27_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave27 scb_axis_mon scb_axis_mon (.*, .model_id(8'd27));
`endif
`ifdef ATCBMC300_SLV28_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave28 scb_axis_mon scb_axis_mon (.*, .model_id(8'd28));
`endif
`ifdef ATCBMC300_SLV29_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave29 scb_axis_mon scb_axis_mon (.*, .model_id(8'd29));
`endif
`ifdef ATCBMC300_SLV30_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave30 scb_axis_mon scb_axis_mon (.*, .model_id(8'd30));
`endif
`ifdef ATCBMC300_SLV31_SUPPORT
bind axi_slave_model : `NDS_SYSTEM.axi_slave31 scb_axis_mon scb_axis_mon (.*, .model_id(8'd31));
`endif
`endif // NDS_SCOREBOARD_EN
// VPERL_GENERATED_END
